.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* NGSPICE file created from tempsensor_rcx.ext - technology: sky130A

.subckt tempsensor_rcx vdd vbe1_out ena vbg vbe2_out vss
X0 a_1429_n4304.t2 a_1429_n4304.t1 vss vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X1 a_495_638.t1 a_495_638.t0 vss vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X2 a_764_n1158.t0 ena.t0 vss.t33 vss.t32 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X3 a_1660_n393# ena.t1 vss vss sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_495_638.t0 XQ_BR1.Emitter.t6 a_1537_2302# vss.t38 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X5 vss a_1660_n393# XQ_BR1.Emitter.t4 vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X6 a_2471_n2640.t1 vbe1_out.t0 vbe1_out.t1 vss.t39 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X7 vss.t35 vss.t34 XQ_BR1.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=19848076,36944
D0 vss.t4 vbe2_out.t3 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X8 a_1537_2302# vbe2_out.t1 vbe2_out.t2 vss.t40 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X9 vss a_1660_n393# x2.input.t0 vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X10 vss a_1660_n393# XQ_BR1.Emitter.t3 vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X11 a_1429_n4304.t0 x2.input.t2 a_2471_n2640.t0 vss.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X12 vss a_1660_n393# XQ_BR1.Emitter.t2 vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
D1 vss.t41 vbg.t0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
D2 vss.t25 vbe1_out.t3 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X13 vss.t24 ena.t2 a_1537_2302# vss.t23 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X14 vss a_1660_n393# XQ_BR1.Emitter.t1 vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X15 vss a_495_638.t0 vbe2_out.t0 vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X16 vss a_506_n1158.t1 a_506_n1158.t2 vss sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X17 vss a_1660_n393# XQ_BR1.Emitter.t0 vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X18 a_1660_n393# a_1660_n393# a_764_n1158.t2 vss.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
D3 vss.t6 ena.t3 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X19 a_1660_n393# a_506_n1158.t3 vss vss sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X20 a_764_n1158.t1 vbg.t1 a_506_n1158.t0 vss.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X21 vss.t37 vss.t36 x2.input.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720 d=19848076,36944
X22 vss.t29 ena.t4 a_2471_n2640.t0 vss.t28 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
X23 vss a_1429_n4304.t1 vbe1_out.t2 vss sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
R0 a_1429_n4304.t2 a_1429_n4304.t1 228.215
R1 a_1429_n4304.t1 a_1429_n4304.t0 85.8993
R2 vss.n126 vss.n125 1.39509e+06
R3 vss.n126 vss.n76 993664
R4 vss.n416 vss.n60 75637.7
R5 vss.n627 vss.n8 33184.6
R6 vss.n49 vss.n35 9483.78
R7 vss.n125 vss.n7 8818.62
R8 vss.n628 vss.n627 8694.85
R9 vss.n125 vss.n35 8027.75
R10 vss.n62 vss.n61 8013.27
R11 vss.n574 vss.n61 8013.27
R12 vss.n572 vss.n62 8013.27
R13 vss.n574 vss.n572 8013.27
R14 vss.n184 vss.n81 8013.27
R15 vss.n556 vss.n81 8013.27
R16 vss.n184 vss.n82 8013.27
R17 vss.n556 vss.n82 8013.27
R18 vss.n414 vss.n179 8013.27
R19 vss.n414 vss.n180 8013.27
R20 vss.n570 vss.n65 8013.27
R21 vss.n570 vss.n66 8013.27
R22 vss.n618 vss.n19 8013.27
R23 vss.n19 vss.n17 8013.27
R24 vss.n18 vss.n17 8013.27
R25 vss.n618 vss.n18 8013.27
R26 vss.n625 vss.n9 8013.27
R27 vss.n625 vss.n10 8013.27
R28 vss.n32 vss.n30 8013.27
R29 vss.n32 vss.n31 8013.27
R30 vss.n628 vss.n7 7452.73
R31 vss.n602 vss.n35 6644.9
R32 vss.n179 vss.n70 6622.68
R33 vss.n70 vss.n65 6622.68
R34 vss.n180 vss.n71 6622.68
R35 vss.n71 vss.n66 6622.68
R36 vss.n14 vss.n9 6622.68
R37 vss.n30 vss.n14 6622.68
R38 vss.n15 vss.n10 6622.68
R39 vss.n31 vss.n15 6622.68
R40 vss.n603 vss.n602 6301.58
R41 vss.n602 vss.n601 6293.61
R42 vss.n629 vss.n628 5221.33
R43 vss.t37 vss.n76 5215.79
R44 vss.n626 vss.t38 2854.26
R45 vss.n594 vss.n37 2798.56
R46 vss.n600 vss.n37 2798.56
R47 vss.n594 vss.n38 2798.56
R48 vss.n600 vss.n38 2798.56
R49 vss.n129 vss.n128 2798.56
R50 vss.n131 vss.n129 2798.56
R51 vss.n132 vss.n128 2798.56
R52 vss.n132 vss.n131 2798.56
R53 vss.n412 vss.n182 2713.02
R54 vss.n619 vss.n16 2681.95
R55 vss.t23 vss.t40 2681.95
R56 vss.n33 vss.n29 2681.95
R57 vss.t37 vss.t39 2318.31
R58 vss.n528 vss.n94 1548.43
R59 vss.n302 vss.n93 1471.78
R60 vss.n248 vss.n247 1450.55
R61 vss.n247 vss.n246 1450.55
R62 vss.n246 vss.n234 1450.55
R63 vss.n240 vss.n234 1450.55
R64 vss.n611 vss.n27 1407.97
R65 vss.n611 vss.n28 1407.97
R66 vss.n610 vss.n27 1407.97
R67 vss.n610 vss.n28 1407.97
R68 vss.n578 vss.n58 1407.97
R69 vss.n578 vss.n59 1407.97
R70 vss.n579 vss.n58 1407.97
R71 vss.n579 vss.n59 1407.97
R72 vss.n585 vss.n51 1407.97
R73 vss.n585 vss.n52 1407.97
R74 vss.n51 vss.n50 1407.97
R75 vss.n52 vss.n50 1407.97
R76 vss.n587 vss.n44 1407.97
R77 vss.n591 vss.n44 1407.97
R78 vss.n587 vss.n45 1407.97
R79 vss.n591 vss.n45 1407.97
R80 vss.n620 vss.n14 1390.59
R81 vss.n620 vss.n15 1390.59
R82 vss.n564 vss.n70 1390.59
R83 vss.n564 vss.n71 1390.59
R84 vss.n522 vss.n94 1379.79
R85 vss.n522 vss.n521 1379.79
R86 vss.n521 vss.n520 1379.79
R87 vss.n520 vss.n99 1379.79
R88 vss.n631 vss.n5 1379.79
R89 vss.n631 vss.n630 1379.79
R90 vss.n303 vss.n6 1379.79
R91 vss.n303 vss.n302 1379.79
R92 vss.n529 vss.n93 1211.15
R93 vss.n529 vss.n528 1195.82
R94 vss.n240 vss.n239 1144.93
R95 vss.n630 vss.n629 1042.51
R96 vss.n608 vss.n26 1028.14
R97 vss.t32 vss.n64 899.119
R98 vss.n124 vss.n80 883.88
R99 vss.n183 vss.t29 872.783
R100 vss.n22 vss.t24 872.783
R101 vss.n605 vss.n26 806.4
R102 vss.n183 vss.n69 791.34
R103 vss.n22 vss.n13 791.34
R104 vss.n99 vss.n0 804.317
R105 vss.n253 vss.n252 760.077
R106 vss.n253 vss.n227 760.077
R107 vss.n374 vss.n227 760.077
R108 vss.n375 vss.n374 760.077
R109 vss.n376 vss.n375 760.077
R110 vss.n376 vss.n209 760.077
R111 vss.n389 vss.n210 760.077
R112 vss.n217 vss.n210 760.077
R113 vss.n217 vss.n177 760.077
R114 vss.n418 vss.n177 760.077
R115 vss.n418 vss.n417 760.077
R116 vss.n239 vss.n238 733.638
R117 vss.t35 vss.n5 720.558
R118 vss.n252 vss.n8 709.405
R119 vss.n559 vss.n558 609.442
R120 vss.n397 vss.n89 602.201
R121 vss.n90 vss.n89 599.201
R122 vss.n568 vss.n567 596.898
R123 vss.n517 vss.n100 585
R124 vss.n100 vss.n99 585
R125 vss.n519 vss.n518 585
R126 vss.n520 vss.n519 585
R127 vss.n101 vss.n98 585
R128 vss.n521 vss.n98 585
R129 vss.n523 vss.n97 585
R130 vss.n523 vss.n522 585
R131 vss.n110 vss.n103 585
R132 vss.n508 vss.n105 585
R133 vss.n510 vss.n509 585
R134 vss.n512 vss.n104 585
R135 vss.n513 vss.n102 585
R136 vss.n516 vss.n515 585
R137 vss.n505 vss.n504 585
R138 vss.n148 vss.n75 585
R139 vss.n147 vss.n144 585
R140 vss.n479 vss.n478 585
R141 vss.n482 vss.n481 585
R142 vss.n142 vss.n139 585
R143 vss.n136 vss.n122 585
R144 vss.n490 vss.n489 585
R145 vss.n493 vss.n492 585
R146 vss.n121 vss.n118 585
R147 vss.n115 vss.n111 585
R148 vss.n501 vss.n500 585
R149 vss.n501 vss.n80 585
R150 vss.n502 vss.n109 585
R151 vss.n562 vss.n561 585
R152 vss.n549 vss.n73 585
R153 vss.n73 vss.n72 585
R154 vss.n548 vss.n547 585
R155 vss.n547 vss.n546 585
R156 vss.n544 vss.n83 585
R157 vss.n545 vss.n544 585
R158 vss.n543 vss.n542 585
R159 vss.n543 vss.n78 585
R160 vss.n541 vss.n84 585
R161 vss.n84 vss.n79 585
R162 vss.n540 vss.n539 585
R163 vss.n539 vss.n538 585
R164 vss.n86 vss.n85 585
R165 vss.n537 vss.n86 585
R166 vss.n535 vss.n534 585
R167 vss.n536 vss.n535 585
R168 vss.n533 vss.n88 585
R169 vss.n88 vss.n87 585
R170 vss.n249 vss.n233 585
R171 vss.n249 vss.n248 585
R172 vss.n251 vss.n231 585
R173 vss.n252 vss.n251 585
R174 vss.n255 vss.n254 585
R175 vss.n254 vss.n253 585
R176 vss.n229 vss.n228 585
R177 vss.n228 vss.n227 585
R178 vss.n373 vss.n372 585
R179 vss.n374 vss.n373 585
R180 vss.n226 vss.n225 585
R181 vss.n375 vss.n226 585
R182 vss.n378 vss.n377 585
R183 vss.n377 vss.n376 585
R184 vss.n222 vss.n211 585
R185 vss.n211 vss.n209 585
R186 vss.n388 vss.n387 585
R187 vss.n389 vss.n388 585
R188 vss.n214 vss.n212 585
R189 vss.n212 vss.n210 585
R190 vss.n219 vss.n218 585
R191 vss.n218 vss.n217 585
R192 vss.n175 vss.n173 585
R193 vss.n177 vss.n175 585
R194 vss.n420 vss.n419 585
R195 vss.n419 vss.n418 585
R196 vss.n181 vss.n176 585
R197 vss.n417 vss.n176 585
R198 vss.n242 vss.n241 585
R199 vss.n241 vss.n240 585
R200 vss.n243 vss.n235 585
R201 vss.n235 vss.n234 585
R202 vss.n245 vss.n244 585
R203 vss.n246 vss.n245 585
R204 vss.n236 vss.n232 585
R205 vss.n247 vss.n232 585
R206 vss.n525 vss.n524 585
R207 vss.n524 vss.n94 585
R208 vss.n398 vss.n392 585
R209 vss.n399 vss.n398 585
R210 vss.n402 vss.n401 585
R211 vss.n401 vss.n400 585
R212 vss.n403 vss.n391 585
R213 vss.n391 vss.n390 585
R214 vss.n405 vss.n404 585
R215 vss.n406 vss.n405 585
R216 vss.n193 vss.n191 585
R217 vss.n407 vss.n193 585
R218 vss.n410 vss.n409 585
R219 vss.n409 vss.n408 585
R220 vss.n192 vss.n190 585
R221 vss.n208 vss.n192 585
R222 vss.n206 vss.n205 585
R223 vss.n207 vss.n206 585
R224 vss.n204 vss.n195 585
R225 vss.n195 vss.n194 585
R226 vss.n203 vss.n202 585
R227 vss.n202 vss.n201 585
R228 vss.n199 vss.n196 585
R229 vss.n200 vss.n199 585
R230 vss.n198 vss.n197 585
R231 vss.n198 vss.n178 585
R232 vss.n532 vss.n531 585
R233 vss.n531 vss.n530 585
R234 vss.n395 vss.n394 585
R235 vss.n454 vss.n158 585
R236 vss.n450 vss.n449 585
R237 vss.n447 vss.n446 585
R238 vss.n284 vss.n279 585
R239 vss.n278 vss.n276 585
R240 vss.n297 vss.n271 585
R241 vss.n343 vss.n267 585
R242 vss.n310 vss.n263 585
R243 vss.n311 vss.n262 585
R244 vss.n336 vss.n313 585
R245 vss.n337 vss.n336 585
R246 vss.n339 vss.n262 585
R247 vss.n340 vss.n263 585
R248 vss.n343 vss.n342 585
R249 vss.n298 vss.n297 585
R250 vss.n281 vss.n276 585
R251 vss.n284 vss.n283 585
R252 vss.n446 vss.n162 585
R253 vss.n451 vss.n450 585
R254 vss.n454 vss.n453 585
R255 vss.n394 vss.n161 585
R256 vss.n306 vss.n299 585
R257 vss.n302 vss.n299 585
R258 vss.n305 vss.n304 585
R259 vss.n304 vss.n303 585
R260 vss.n301 vss.n300 585
R261 vss.n301 vss.n6 585
R262 vss.n4 vss.n2 585
R263 vss.n630 vss.n4 585
R264 vss.n633 vss.n632 585
R265 vss.n632 vss.n631 585
R266 vss.n3 vss.n1 585
R267 vss.n5 vss.n3 585
R268 vss.n238 vss.n237 585
R269 vss.n308 vss.n307 585
R270 vss.n308 vss.n93 585
R271 vss.n527 vss.n526 585
R272 vss.n528 vss.n527 585
R273 vss.n627 vss.n626 551.874
R274 vss.n584 vss.n53 533.208
R275 vss.n413 vss.n68 520.659
R276 vss.n624 vss.n623 520.659
R277 vss.t35 vss.n389 515.163
R278 vss.n607 vss.n12 437.159
R279 vss.n416 vss.n415 427.812
R280 vss.n530 vss.n529 427.812
R281 vss.n567 vss.n566 411.483
R282 vss.n622 vss.n12 411.483
R283 vss.n566 vss.n68 409.976
R284 vss.n623 vss.n622 409.976
R285 vss.n248 vss.n8 386.813
R286 vss.t32 vss.n571 354.661
R287 vss.n239 vss.t35 337.858
R288 vss.n629 vss.n6 337.283
R289 vss.n529 vss.n92 336.171
R290 vss.n529 vss.n77 331.916
R291 vss.t37 vss.n77 327.661
R292 vss.t4 vss.n34 324.632
R293 vss.t35 vss.n92 323.404
R294 vss.t4 vss.n603 322.135
R295 vss.n50 vss.n46 311.077
R296 vss.n592 vss.n43 304.786
R297 vss.n103 vss.n0 250.21
R298 vss.n34 vss.n33 297.163
R299 vss.n603 vss.n28 294.998
R300 vss.n591 vss.n590 292.5
R301 vss.n592 vss.n591 292.5
R302 vss.n589 vss.n45 292.5
R303 vss.t25 vss.n45 292.5
R304 vss.n588 vss.n587 292.5
R305 vss.n587 vss.n586 292.5
R306 vss.n47 vss.n44 292.5
R307 vss.t25 vss.n44 292.5
R308 vss.n582 vss.n52 292.5
R309 vss.n52 vss.n42 292.5
R310 vss.t6 vss.n50 292.5
R311 vss.n54 vss.n51 292.5
R312 vss.n51 vss.n48 292.5
R313 vss.n585 vss.n584 292.5
R314 vss.t6 vss.n585 292.5
R315 vss.n59 vss.n57 292.5
R316 vss.n59 vss.n36 292.5
R317 vss.n580 vss.n579 292.5
R318 vss.n579 vss.t41 292.5
R319 vss.n58 vss.n56 292.5
R320 vss.n58 vss.n43 292.5
R321 vss.n578 vss.n577 292.5
R322 vss.t41 vss.n578 292.5
R323 vss.n608 vss.n28 292.5
R324 vss.n610 vss.n609 292.5
R325 vss.t4 vss.n610 292.5
R326 vss.n606 vss.n27 292.5
R327 vss.n34 vss.n27 292.5
R328 vss.n612 vss.n611 292.5
R329 vss.n611 vss.t4 292.5
R330 vss.n605 vss.n604 288
R331 vss.n503 vss.n80 263.904
R332 vss.n476 vss.n475 258.334
R333 vss.n441 vss.n440 258.334
R334 vss.n531 vss.n90 257.466
R335 vss.n198 vss.n176 257.466
R336 vss.n506 vss.n108 254.34
R337 vss.n107 vss.n103 254.34
R338 vss.n511 vss.n103 254.34
R339 vss.n514 vss.n103 254.34
R340 vss.n143 vss.n80 254.34
R341 vss.n480 vss.n80 254.34
R342 vss.n141 vss.n80 254.34
R343 vss.n491 vss.n80 254.34
R344 vss.n120 vss.n80 254.34
R345 vss.n560 vss.n74 254.34
R346 vss.n396 vss.n92 254.34
R347 vss.n448 vss.n92 254.34
R348 vss.n164 vss.n92 254.34
R349 vss.n277 vss.n92 254.34
R350 vss.n309 vss.n92 254.34
R351 vss.n312 vss.n92 254.34
R352 vss.n338 vss.n77 254.34
R353 vss.n341 vss.n77 254.34
R354 vss.n269 vss.n77 254.34
R355 vss.n282 vss.n77 254.34
R356 vss.n452 vss.n77 254.34
R357 vss.n160 vss.n77 254.34
R358 vss.n559 vss.n75 251.614
R359 vss.n398 vss.n397 251.614
R360 vss.n415 vss.n178 250.952
R361 vss.n459 vss.n458 250
R362 vss.n126 vss.t10 249.37
R363 vss.t35 vss.n209 244.915
R364 vss.n557 vss.n64 234.131
R365 vss.n200 vss.n178 215.101
R366 vss.n201 vss.n200 215.101
R367 vss.n201 vss.n194 215.101
R368 vss.n207 vss.n194 215.101
R369 vss.n208 vss.n207 215.101
R370 vss.n408 vss.n407 215.101
R371 vss.n407 vss.n406 215.101
R372 vss.n406 vss.n390 215.101
R373 vss.n400 vss.n390 215.101
R374 vss.n400 vss.n399 215.101
R375 vss.n530 vss.n87 215.101
R376 vss.n536 vss.n87 215.101
R377 vss.n537 vss.n536 215.101
R378 vss.n538 vss.n537 215.101
R379 vss.n538 vss.n79 215.101
R380 vss.n545 vss.n78 215.101
R381 vss.n546 vss.n545 215.101
R382 vss.n546 vss.n72 215.101
R383 vss.n615 vss.n24 212.103
R384 vss.n524 vss.n95 195.049
R385 vss.n250 vss.n249 195.049
R386 vss.n617 vss.n616 194.21
R387 vss.n554 vss.n553 192.385
R388 vss.n504 vss.n110 187.249
R389 vss.n308 vss.n299 187.249
R390 vss.n320 vss.n319 185
R391 vss.n322 vss.n321 185
R392 vss.n324 vss.n318 185
R393 vss.n326 vss.n325 185
R394 vss.n327 vss.n316 185
R395 vss.n329 vss.n328 185
R396 vss.n331 vss.n315 185
R397 vss.n332 vss.n314 185
R398 vss.n332 vss.t36 185
R399 vss.n334 vss.n333 185
R400 vss.n475 vss.n150 185
R401 vss.n473 vss.n472 185
R402 vss.n471 vss.n151 185
R403 vss.n470 vss.n469 185
R404 vss.n467 vss.n152 185
R405 vss.n465 vss.n464 185
R406 vss.n463 vss.n153 185
R407 vss.n462 vss.n461 185
R408 vss.n459 vss.n154 185
R409 vss.n459 vss.t36 185
R410 vss.n477 vss.n476 185
R411 vss.n140 vss.n138 185
R412 vss.n484 vss.n483 185
R413 vss.n486 vss.n137 185
R414 vss.n488 vss.n487 185
R415 vss.n119 vss.n117 185
R416 vss.n495 vss.n494 185
R417 vss.n497 vss.n116 185
R418 vss.n499 vss.n498 185
R419 vss.n440 vss.n167 185
R420 vss.n438 vss.n437 185
R421 vss.n436 vss.n168 185
R422 vss.n435 vss.n434 185
R423 vss.n432 vss.n169 185
R424 vss.n430 vss.n429 185
R425 vss.n428 vss.n170 185
R426 vss.n427 vss.n426 185
R427 vss.n424 vss.n171 185
R428 vss.n351 vss.n260 185
R429 vss.n353 vss.n352 185
R430 vss.n355 vss.n354 185
R431 vss.n358 vss.n357 185
R432 vss.n359 vss.n258 185
R433 vss.n361 vss.n360 185
R434 vss.n363 vss.n257 185
R435 vss.n365 vss.n364 185
R436 vss.n367 vss.n366 185
R437 vss.n370 vss.n369 185
R438 vss.n371 vss.n224 185
R439 vss.n380 vss.n379 185
R440 vss.n382 vss.n223 185
R441 vss.n383 vss.n213 185
R442 vss.n386 vss.n385 185
R443 vss.n221 vss.n220 185
R444 vss.n216 vss.n172 185
R445 vss.n422 vss.n421 185
R446 vss.n441 vss.n159 185
R447 vss.n443 vss.n157 185
R448 vss.n445 vss.n444 185
R449 vss.n280 vss.n275 185
R450 vss.n293 vss.n292 185
R451 vss.n296 vss.n295 185
R452 vss.n274 vss.n268 185
R453 vss.n266 vss.n261 185
R454 vss.n349 vss.n348 185
R455 vss.n347 vss.n346 185
R456 vss.n345 vss.n344 185
R457 vss.n287 vss.n270 185
R458 vss.n288 vss.n272 185
R459 vss.n291 vss.n290 185
R460 vss.n286 vss.n165 185
R461 vss.n163 vss.n156 185
R462 vss.n456 vss.n455 185
R463 vss.n458 vss.n155 185
R464 vss.n502 vss.n501 175.546
R465 vss.n501 vss.n111 175.546
R466 vss.n492 vss.n121 175.546
R467 vss.n490 vss.n122 175.546
R468 vss.n481 vss.n142 175.546
R469 vss.n479 vss.n144 175.546
R470 vss.n531 vss.n88 175.546
R471 vss.n535 vss.n88 175.546
R472 vss.n535 vss.n86 175.546
R473 vss.n539 vss.n86 175.546
R474 vss.n539 vss.n84 175.546
R475 vss.n543 vss.n84 175.546
R476 vss.n544 vss.n543 175.546
R477 vss.n547 vss.n544 175.546
R478 vss.n547 vss.n73 175.546
R479 vss.n561 vss.n73 175.546
R480 vss.n340 vss.n339 175.546
R481 vss.n342 vss.n298 175.546
R482 vss.n283 vss.n281 175.546
R483 vss.n451 vss.n162 175.546
R484 vss.n453 vss.n161 175.546
R485 vss.n524 vss.n523 175.546
R486 vss.n523 vss.n98 175.546
R487 vss.n519 vss.n98 175.546
R488 vss.n519 vss.n100 175.546
R489 vss.n515 vss.n100 175.546
R490 vss.n513 vss.n512 175.546
R491 vss.n510 vss.n105 175.546
R492 vss.n311 vss.n310 175.546
R493 vss.n271 vss.n267 175.546
R494 vss.n279 vss.n278 175.546
R495 vss.n449 vss.n447 175.546
R496 vss.n395 vss.n158 175.546
R497 vss.n199 vss.n198 175.546
R498 vss.n202 vss.n199 175.546
R499 vss.n202 vss.n195 175.546
R500 vss.n206 vss.n195 175.546
R501 vss.n206 vss.n192 175.546
R502 vss.n409 vss.n192 175.546
R503 vss.n409 vss.n193 175.546
R504 vss.n405 vss.n193 175.546
R505 vss.n405 vss.n391 175.546
R506 vss.n401 vss.n391 175.546
R507 vss.n401 vss.n398 175.546
R508 vss.n254 vss.n228 175.546
R509 vss.n373 vss.n228 175.546
R510 vss.n373 vss.n226 175.546
R511 vss.n377 vss.n226 175.546
R512 vss.n377 vss.n211 175.546
R513 vss.n388 vss.n211 175.546
R514 vss.n388 vss.n212 175.546
R515 vss.n218 vss.n212 175.546
R516 vss.n218 vss.n175 175.546
R517 vss.n419 vss.n175 175.546
R518 vss.n419 vss.n176 175.546
R519 vss.n249 vss.n232 175.546
R520 vss.n245 vss.n232 175.546
R521 vss.n245 vss.n235 175.546
R522 vss.n241 vss.n235 175.546
R523 vss.n241 vss.n238 175.546
R524 vss.n238 vss.n3 175.546
R525 vss.n632 vss.n3 175.546
R526 vss.n632 vss.n4 175.546
R527 vss.n301 vss.n4 175.546
R528 vss.n304 vss.n301 175.546
R529 vss.n304 vss.n299 175.546
R530 vss.n581 vss.n55 172.405
R531 vss.n16 vss.t38 172.304
R532 vss.n619 vss.t23 172.304
R533 vss.n29 vss.t40 172.304
R534 vss.t5 vss.n91 164.911
R535 vss.n369 vss.n367 163.333
R536 vss.t41 vss.t9 153.779
R537 vss.n108 vss.n107 152.643
R538 vss.n563 vss.n562 150.571
R539 vss.n346 vss.n345 150
R540 vss.n288 vss.n287 150
R541 vss.n290 vss.n286 150
R542 vss.n456 vss.n156 150
R543 vss.n333 vss.n332 150
R544 vss.n332 vss.n331 150
R545 vss.n329 vss.n316 150
R546 vss.n325 vss.n324 150
R547 vss.n322 vss.n319 150
R548 vss.n498 vss.n497 150
R549 vss.n495 vss.n117 150
R550 vss.n487 vss.n486 150
R551 vss.n484 vss.n138 150
R552 vss.n461 vss.n459 150
R553 vss.n465 vss.n153 150
R554 vss.n469 vss.n467 150
R555 vss.n473 vss.n151 150
R556 vss.n349 vss.n261 150
R557 vss.n295 vss.n274 150
R558 vss.n293 vss.n275 150
R559 vss.n444 vss.n443 150
R560 vss.n426 vss.n424 150
R561 vss.n430 vss.n170 150
R562 vss.n434 vss.n432 150
R563 vss.n438 vss.n168 150
R564 vss.n380 vss.n224 150
R565 vss.n383 vss.n382 150
R566 vss.n385 vss.n221 150
R567 vss.n422 vss.n172 150
R568 vss.n364 vss.n363 150
R569 vss.n361 vss.n258 150
R570 vss.n357 vss.n355 150
R571 vss.n352 vss.n351 150
R572 vss.n617 vss.n22 147.888
R573 vss.n529 vss.n91 138.62
R574 vss.n586 vss.n48 138.54
R575 vss.n53 vss.n46 136.534
R576 vss.n593 vss.n42 132.998
R577 vss.n313 vss.n308 126.782
R578 vss.n337 vss.n95 124.832
R579 vss.n254 vss.n250 124.832
R580 vss.t41 vss.n60 119.144
R581 vss.n570 vss.n569 117.001
R582 vss.n571 vss.n570 117.001
R583 vss.n556 vss.n555 117.001
R584 vss.n557 vss.n556 117.001
R585 vss.n575 vss.n574 117.001
R586 vss.n574 vss.n573 117.001
R587 vss.n145 vss.n62 117.001
R588 vss.n124 vss.n62 117.001
R589 vss.n131 vss.n130 117.001
R590 vss.n131 vss.n64 117.001
R591 vss.n133 vss.n132 117.001
R592 vss.n132 vss.t10 117.001
R593 vss.n128 vss.n113 117.001
R594 vss.n128 vss.n127 117.001
R595 vss.n129 vss.n106 117.001
R596 vss.n129 vss.t10 117.001
R597 vss.n600 vss.n599 117.001
R598 vss.n601 vss.n600 117.001
R599 vss.n597 vss.n38 117.001
R600 vss.t9 vss.n38 117.001
R601 vss.n595 vss.n594 117.001
R602 vss.n594 vss.n593 117.001
R603 vss.n39 vss.n37 117.001
R604 vss.t9 vss.n37 117.001
R605 vss.n565 vss.n564 117.001
R606 vss.n564 vss.n563 117.001
R607 vss.n414 vss.n413 117.001
R608 vss.n415 vss.n414 117.001
R609 vss.n185 vss.n184 117.001
R610 vss.n184 vss.n91 117.001
R611 vss.n21 vss.n18 117.001
R612 vss.n18 vss.n16 117.001
R613 vss.n625 vss.n624 117.001
R614 vss.n626 vss.n625 117.001
R615 vss.n621 vss.n620 117.001
R616 vss.n620 vss.n619 117.001
R617 vss.n616 vss.n19 117.001
R618 vss.n29 vss.n19 117.001
R619 vss.n32 vss.n25 117.001
R620 vss.n33 vss.n32 117.001
R621 vss.n49 vss.t25 114.987
R622 vss.n399 vss.t5 114.721
R623 vss.n54 vss.n53 114.162
R624 vss.n408 vss.t35 112.331
R625 vss.t37 vss.n78 112.331
R626 vss.t37 vss.n80 105.29
R627 vss.n599 vss.n39 104.534
R628 vss.t35 vss.n208 102.77
R629 vss.t37 vss.n79 102.77
R630 vss.t39 vss.n557 95.5924
R631 vss.n609 vss.n608 91.4829
R632 vss.n589 vss.n588 91.4829
R633 vss.n580 vss.n57 91.4829
R634 vss.n624 vss.n11 89.8066
R635 vss.n127 vss.n126 87.2801
R636 vss.n507 vss.n106 85.6701
R637 vss.n123 vss.n106 82.824
R638 vss.n568 vss.n53 82.3356
R639 vss.n413 vss.n412 79.8123
R640 vss.n596 vss.n39 79.8123
R641 vss.n40 vss.t33 79.2195
R642 vss.n120 vss.n111 76.3222
R643 vss.n492 vss.n491 76.3222
R644 vss.n141 vss.n122 76.3222
R645 vss.n481 vss.n480 76.3222
R646 vss.n144 vss.n143 76.3222
R647 vss.n560 vss.n559 76.3222
R648 vss.n338 vss.n337 76.3222
R649 vss.n341 vss.n340 76.3222
R650 vss.n298 vss.n269 76.3222
R651 vss.n283 vss.n282 76.3222
R652 vss.n452 vss.n451 76.3222
R653 vss.n161 vss.n160 76.3222
R654 vss.n514 vss.n513 76.3222
R655 vss.n511 vss.n510 76.3222
R656 vss.n110 vss.n108 76.3222
R657 vss.n107 vss.n105 76.3222
R658 vss.n512 vss.n511 76.3222
R659 vss.n515 vss.n514 76.3222
R660 vss.n143 vss.n75 76.3222
R661 vss.n480 vss.n479 76.3222
R662 vss.n142 vss.n141 76.3222
R663 vss.n491 vss.n490 76.3222
R664 vss.n121 vss.n120 76.3222
R665 vss.n561 vss.n560 76.3222
R666 vss.n312 vss.n311 76.3222
R667 vss.n309 vss.n267 76.3222
R668 vss.n278 vss.n277 76.3222
R669 vss.n447 vss.n164 76.3222
R670 vss.n448 vss.n158 76.3222
R671 vss.n397 vss.n396 76.3222
R672 vss.n396 vss.n395 76.3222
R673 vss.n449 vss.n448 76.3222
R674 vss.n279 vss.n164 76.3222
R675 vss.n277 vss.n271 76.3222
R676 vss.n310 vss.n309 76.3222
R677 vss.n313 vss.n312 76.3222
R678 vss.n339 vss.n338 76.3222
R679 vss.n342 vss.n341 76.3222
R680 vss.n281 vss.n269 76.3222
R681 vss.n282 vss.n162 76.3222
R682 vss.n453 vss.n452 76.3222
R683 vss.n160 vss.n90 76.3222
R684 vss.n423 vss.n422 74.5978
R685 vss.n424 vss.n423 74.5978
R686 vss.n558 vss.t28 73.6705
R687 vss.n569 vss.n67 72.6492
R688 vss.n565 vss.n69 70.4005
R689 vss.n621 vss.n13 70.4005
R690 vss.n498 vss.n114 69.3109
R691 vss.n319 vss.n114 69.3109
R692 vss.n350 vss.n349 69.3109
R693 vss.n351 vss.n350 69.3109
R694 vss.n571 vss.n48 67.8846
R695 vss.n323 vss.t36 65.8183
R696 vss.n317 vss.t36 65.8183
R697 vss.n330 vss.t36 65.8183
R698 vss.n474 vss.t36 65.8183
R699 vss.n468 vss.t36 65.8183
R700 vss.n466 vss.t36 65.8183
R701 vss.n460 vss.t36 65.8183
R702 vss.n146 vss.t36 65.8183
R703 vss.n485 vss.t36 65.8183
R704 vss.n135 vss.t36 65.8183
R705 vss.n496 vss.t36 65.8183
R706 vss.n439 vss.t34 65.8183
R707 vss.n433 vss.t34 65.8183
R708 vss.n431 vss.t34 65.8183
R709 vss.n425 vss.t34 65.8183
R710 vss.n259 vss.t34 65.8183
R711 vss.n356 vss.t34 65.8183
R712 vss.n362 vss.t34 65.8183
R713 vss.n230 vss.t34 65.8183
R714 vss.n368 vss.t34 65.8183
R715 vss.n381 vss.t34 65.8183
R716 vss.n384 vss.t34 65.8183
R717 vss.n215 vss.t34 65.8183
R718 vss.n442 vss.t34 65.8183
R719 vss.t34 vss.n166 65.8183
R720 vss.n294 vss.t34 65.8183
R721 vss.n273 vss.t34 65.8183
R722 vss.n265 vss.t36 65.8183
R723 vss.n289 vss.t36 65.8183
R724 vss.n285 vss.t36 65.8183
R725 vss.n457 vss.t36 65.8183
R726 vss.n55 vss.n54 64.6924
R727 vss.n563 vss.n72 64.5307
R728 vss.n264 vss.t36 64.1729
R729 vss.n573 vss.n60 58.1869
R730 vss.t36 vss.n114 57.8461
R731 vss.n350 vss.t34 57.8461
R732 vss.n504 vss.n503 57.1945
R733 vss.n503 vss.n502 57.1945
R734 vss.n346 vss.n264 56.6572
R735 vss.n333 vss.n264 56.6572
R736 vss.n423 vss.t34 55.2026
R737 vss.n345 vss.n265 53.3664
R738 vss.n289 vss.n288 53.3664
R739 vss.n286 vss.n285 53.3664
R740 vss.n457 vss.n456 53.3664
R741 vss.n330 vss.n329 53.3664
R742 vss.n325 vss.n317 53.3664
R743 vss.n323 vss.n322 53.3664
R744 vss.n324 vss.n323 53.3664
R745 vss.n317 vss.n316 53.3664
R746 vss.n331 vss.n330 53.3664
R747 vss.n496 vss.n495 53.3664
R748 vss.n487 vss.n135 53.3664
R749 vss.n485 vss.n484 53.3664
R750 vss.n476 vss.n146 53.3664
R751 vss.n460 vss.n153 53.3664
R752 vss.n466 vss.n465 53.3664
R753 vss.n468 vss.n151 53.3664
R754 vss.n474 vss.n473 53.3664
R755 vss.n475 vss.n474 53.3664
R756 vss.n469 vss.n468 53.3664
R757 vss.n467 vss.n466 53.3664
R758 vss.n461 vss.n460 53.3664
R759 vss.n146 vss.n138 53.3664
R760 vss.n486 vss.n485 53.3664
R761 vss.n135 vss.n117 53.3664
R762 vss.n497 vss.n496 53.3664
R763 vss.n274 vss.n273 53.3664
R764 vss.n294 vss.n293 53.3664
R765 vss.n444 vss.n166 53.3664
R766 vss.n442 vss.n441 53.3664
R767 vss.n426 vss.n425 53.3664
R768 vss.n431 vss.n430 53.3664
R769 vss.n434 vss.n433 53.3664
R770 vss.n439 vss.n438 53.3664
R771 vss.n440 vss.n439 53.3664
R772 vss.n433 vss.n168 53.3664
R773 vss.n432 vss.n431 53.3664
R774 vss.n425 vss.n170 53.3664
R775 vss.n369 vss.n368 53.3664
R776 vss.n381 vss.n380 53.3664
R777 vss.n384 vss.n383 53.3664
R778 vss.n221 vss.n215 53.3664
R779 vss.n367 vss.n230 53.3664
R780 vss.n363 vss.n362 53.3664
R781 vss.n356 vss.n258 53.3664
R782 vss.n355 vss.n259 53.3664
R783 vss.n352 vss.n259 53.3664
R784 vss.n357 vss.n356 53.3664
R785 vss.n362 vss.n361 53.3664
R786 vss.n364 vss.n230 53.3664
R787 vss.n368 vss.n224 53.3664
R788 vss.n382 vss.n381 53.3664
R789 vss.n385 vss.n384 53.3664
R790 vss.n215 vss.n172 53.3664
R791 vss.n443 vss.n442 53.3664
R792 vss.n275 vss.n166 53.3664
R793 vss.n295 vss.n294 53.3664
R794 vss.n273 vss.n261 53.3664
R795 vss.n287 vss.n265 53.3664
R796 vss.n290 vss.n289 53.3664
R797 vss.n285 vss.n156 53.3664
R798 vss.n458 vss.n457 53.3664
R799 vss.n609 vss.n607 52.6144
R800 vss.t37 vss.n0 24.7457
R801 vss.n417 vss.n416 50.6723
R802 vss.n576 vss.n57 48.6907
R803 vss.n590 vss.n589 48.0123
R804 vss.n553 vss.n552 45.8245
R805 vss.n24 vss.n23 45.8245
R806 vss.n599 vss.n598 45.5534
R807 vss.n598 vss.n40 45.4279
R808 vss.n576 vss.n575 44.0476
R809 vss.n581 vss.n580 43.432
R810 vss.n584 vss.n583 42.5417
R811 vss.n588 vss.n47 41.5855
R812 vss.n586 vss.t6 41.5622
R813 vss.t25 vss.n42 41.5622
R814 vss.n590 vss.n46 32.1774
R815 vss.n566 vss.n565 31.557
R816 vss.n622 vss.n621 31.557
R817 vss.n582 vss.n46 28.1851
R818 vss.t9 vss.n43 26.3229
R819 vss.n607 vss.n604 24.3205
R820 vss.n577 vss.n56 24.1034
R821 vss.t6 vss.n49 23.5521
R822 vss.n551 vss.n81 20.6635
R823 vss.n76 vss.n7 20.5966
R824 vss.n567 vss.n66 18.8715
R825 vss.t39 vss.n66 18.8715
R826 vss.n553 vss.n65 18.8715
R827 vss.t39 vss.n65 18.8715
R828 vss.n572 vss.n63 18.8715
R829 vss.n572 vss.t32 18.8715
R830 vss.n61 vss.n41 18.8715
R831 vss.t32 vss.n61 18.8715
R832 vss.n180 vss.n68 18.8715
R833 vss.t5 vss.n180 18.8715
R834 vss.n186 vss.n179 18.8715
R835 vss.t5 vss.n179 18.8715
R836 vss.n552 vss.n82 18.8715
R837 vss.n82 vss.t28 18.8715
R838 vss.n81 vss.t28 18.8715
R839 vss.n618 vss.n617 18.8715
R840 vss.t23 vss.n618 18.8715
R841 vss.n20 vss.n9 18.8715
R842 vss.n9 vss.t38 18.8715
R843 vss.n31 vss.n12 18.8715
R844 vss.n31 vss.t40 18.8715
R845 vss.n623 vss.n10 18.8715
R846 vss.n10 vss.t38 18.8715
R847 vss.n30 vss.n24 18.8715
R848 vss.n30 vss.t40 18.8715
R849 vss.n23 vss.n17 18.8715
R850 vss.t23 vss.n17 18.8715
R851 vss.n47 vss.n46 18.4642
R852 vss.n558 vss.t37 17.5414
R853 vss.n616 vss.n615 17.1248
R854 vss.n613 vss.n25 16.8005
R855 vss.n615 vss.n614 16.2422
R856 vss.n606 vss.n605 16.0716
R857 vss.n334 vss.n314 16.0005
R858 vss.n315 vss.n314 16.0005
R859 vss.n328 vss.n315 16.0005
R860 vss.n328 vss.n327 16.0005
R861 vss.n327 vss.n326 16.0005
R862 vss.n321 vss.n318 16.0005
R863 vss.n321 vss.n320 16.0005
R864 vss.n462 vss.n154 16.0005
R865 vss.n463 vss.n462 16.0005
R866 vss.n464 vss.n463 16.0005
R867 vss.n464 vss.n152 16.0005
R868 vss.n470 vss.n152 16.0005
R869 vss.n471 vss.n470 16.0005
R870 vss.n472 vss.n471 16.0005
R871 vss.n472 vss.n150 16.0005
R872 vss.n427 vss.n171 16.0005
R873 vss.n428 vss.n427 16.0005
R874 vss.n429 vss.n428 16.0005
R875 vss.n429 vss.n169 16.0005
R876 vss.n435 vss.n169 16.0005
R877 vss.n436 vss.n435 16.0005
R878 vss.n437 vss.n436 16.0005
R879 vss.n437 vss.n167 16.0005
R880 vss.n366 vss.n365 16.0005
R881 vss.n365 vss.n257 16.0005
R882 vss.n360 vss.n257 16.0005
R883 vss.n360 vss.n359 16.0005
R884 vss.n359 vss.n358 16.0005
R885 vss.n354 vss.n353 16.0005
R886 vss.n353 vss.n260 16.0005
R887 vss.n562 vss.t28 14.3405
R888 vss.n335 vss.n260 13.5116
R889 vss.n318 vss 12.9783
R890 vss.n320 vss.n112 12.9783
R891 vss.n354 vss 12.9783
R892 vss.n554 vss.n551 12.4625
R893 vss.n101 vss.n97 11.6369
R894 vss.n518 vss.n101 11.6369
R895 vss.n518 vss.n517 11.6369
R896 vss.n517 vss.n516 11.6369
R897 vss.n516 vss.n102 11.6369
R898 vss.n509 vss.n104 11.6369
R899 vss.n509 vss.n508 11.6369
R900 vss.n244 vss.n236 11.6369
R901 vss.n244 vss.n243 11.6369
R902 vss.n243 vss.n242 11.6369
R903 vss.n242 vss.n237 11.6369
R904 vss.n237 vss.n1 11.6369
R905 vss.n633 vss.n2 11.6369
R906 vss.n300 vss.n2 11.6369
R907 vss.n305 vss.n300 11.6369
R908 vss.n508 vss.n507 11.5076
R909 vss.n127 vss.n124 11.0836
R910 vss.n134 vss.n133 10.8757
R911 vss.n133 vss.n123 10.587
R912 vss.n595 vss.n41 10.4978
R913 vss.n104 vss 10.3439
R914 vss vss.n633 10.3439
R915 vss.n130 vss.n41 10.3072
R916 vss.n597 vss.n596 10.202
R917 vss.n555 vss.n63 10.1462
R918 vss.n569 vss.n568 10.0329
R919 vss.n412 vss.n411 10.0283
R920 vss.n393 vss.n154 9.95606
R921 vss.n174 vss.n171 9.77828
R922 vss.n581 vss.n56 9.6005
R923 vss.n598 vss.n597 9.2396
R924 vss.n583 vss.n581 8.8005
R925 vss.n614 vss.n613 8.46733
R926 vss.n189 vss.n186 8.28285
R927 vss.n583 vss.n582 8.0005
R928 vss.n393 vss.n167 7.46717
R929 vss.n614 vss 7.43059
R930 vss.n20 vss.n11 7.34078
R931 vss.n392 vss.n89 7.08135
R932 vss.n150 vss.n149 6.93383
R933 vss.t39 vss.t10 6.92745
R934 vss.n306 vss.n305 6.7857
R935 vss.n532 vss.n89 6.69229
R936 vss.n525 vss.n97 6.08263
R937 vss.n526 vss.n525 5.9581
R938 vss.n307 vss.n306 5.66317
R939 vss.n593 vss.n592 5.54206
R940 vss.n607 vss.n606 5.40494
R941 vss.n307 vss.n96 5.07331
R942 vss.n255 vss.n231 4.64566
R943 vss.n577 vss.n576 4.58811
R944 vss.n526 vss.n96 4.18852
R945 vss.n335 vss.n334 3.91161
R946 vss.n366 vss.n256 3.73383
R947 vss.n372 vss.n370 3.6134
R948 vss.n371 vss.n225 3.6134
R949 vss.n379 vss.n378 3.6134
R950 vss.n223 vss.n222 3.6134
R951 vss.n387 vss.n213 3.6134
R952 vss.n386 vss.n214 3.6134
R953 vss.n220 vss.n219 3.6134
R954 vss.n216 vss.n173 3.6134
R955 vss.n421 vss.n420 3.6134
R956 vss.n197 vss.n196 3.50202
R957 vss.n203 vss.n196 3.50202
R958 vss.n204 vss.n203 3.50202
R959 vss.n205 vss.n204 3.50202
R960 vss.n205 vss.n190 3.50202
R961 vss.n410 vss.n191 3.50202
R962 vss.n404 vss.n191 3.50202
R963 vss.n404 vss.n403 3.50202
R964 vss.n403 vss.n402 3.50202
R965 vss.n402 vss.n392 3.50202
R966 vss.n533 vss.n532 3.4999
R967 vss.n534 vss.n533 3.48086
R968 vss.n534 vss.n85 3.48086
R969 vss.n540 vss.n85 3.48086
R970 vss.n541 vss.n540 3.48086
R971 vss.n542 vss.n541 3.48086
R972 vss.n542 vss.n83 3.48086
R973 vss.n548 vss.n83 3.48086
R974 vss.n549 vss.n548 3.48086
R975 vss.n550 vss.n549 3.44219
R976 vss.n181 vss.n174 3.40695
R977 vss.n552 vss.n69 3.24317
R978 vss.n23 vss.n13 3.24317
R979 vss.n67 vss.n63 3.16329
R980 vss.n613 vss.n612 3.08071
R981 vss.n326 vss 3.02272
R982 vss.n358 vss 3.02272
R983 vss.n256 vss.n229 2.89082
R984 vss.n573 vss.n36 2.77128
R985 vss.n601 vss.n36 2.77128
R986 vss.n411 vss.n410 2.29594
R987 vss.n527 vss.n95 1.951
R988 vss.n251 vss.n250 1.951
R989 vss.n256 vss.n255 1.75534
R990 vss.n182 vss.n181 1.75534
R991 vss.n550 vss.n74 1.74732
R992 vss.n347 vss.n263 1.70392
R993 vss.n344 vss.n343 1.70392
R994 vss.n297 vss.n270 1.70392
R995 vss.n276 vss.n272 1.70392
R996 vss.n291 vss.n284 1.70392
R997 vss.n446 vss.n165 1.70392
R998 vss.n450 vss.n163 1.70392
R999 vss.n455 vss.n454 1.70392
R1000 vss.n394 vss.n155 1.70392
R1001 vss.n197 vss.n182 1.51783
R1002 vss.n335 vss.n262 1.36324
R1003 vss.n505 vss.n109 1.35579
R1004 vss.n118 vss.n116 1.34074
R1005 vss.n494 vss.n493 1.34074
R1006 vss.n489 vss.n119 1.34074
R1007 vss.n139 vss.n137 1.34074
R1008 vss.n483 vss.n482 1.34074
R1009 vss.n478 vss.n140 1.34074
R1010 vss.n188 vss.n187 1.30814
R1011 vss vss.n102 1.29343
R1012 vss vss.n1 1.29343
R1013 vss.n148 vss.n74 1.26544
R1014 vss.n411 vss.n189 1.2497
R1015 vss.n420 vss.n174 1.23921
R1016 vss.n411 vss.n190 1.20658
R1017 vss.n233 vss.n231 1.1876
R1018 vss.n186 vss.n185 1.18125
R1019 vss.n115 vss.n113 1.16003
R1020 vss.n136 vss.n134 1.05462
R1021 vss.n21 vss.n20 1.04695
R1022 vss.n370 vss.n229 1.03276
R1023 vss.n372 vss.n371 1.03276
R1024 vss.n379 vss.n225 1.03276
R1025 vss.n378 vss.n223 1.03276
R1026 vss.n222 vss.n213 1.03276
R1027 vss.n387 vss.n386 1.03276
R1028 vss.n220 vss.n214 1.03276
R1029 vss.n219 vss.n216 1.03276
R1030 vss.n421 vss.n173 1.03276
R1031 vss.n147 vss.n145 1.00944
R1032 vss.n149 vss.n148 0.994382
R1033 vss.n393 vss.n89 0.876546
R1034 vss.n500 vss.n112 0.843794
R1035 vss.n336 vss.n335 0.827876
R1036 vss.n236 vss.n233 0.75019
R1037 vss.n394 vss.n393 0.58453
R1038 vss.n612 vss.n26 0.513869
R1039 vss.n112 vss.n109 0.5125
R1040 vss.n596 vss.n595 0.492808
R1041 vss.n348 vss.n347 0.462857
R1042 vss.n344 vss.n266 0.462857
R1043 vss.n270 vss.n268 0.462857
R1044 vss.n296 vss.n272 0.462857
R1045 vss.n292 vss.n291 0.462857
R1046 vss.n280 vss.n165 0.462857
R1047 vss.n445 vss.n163 0.462857
R1048 vss.n455 vss.n157 0.462857
R1049 vss.n159 vss.n155 0.462857
R1050 vss.n187 vss.n11 0.393952
R1051 vss.n189 vss.n188 0.388
R1052 vss.n130 vss.n123 0.365761
R1053 vss.n149 vss.n147 0.361912
R1054 vss.n506 vss.n505 0.346853
R1055 vss.n551 vss.n550 0.346853
R1056 vss.n477 vss.n145 0.331794
R1057 vss.n185 vss.n183 0.291409
R1058 vss.n488 vss.n134 0.286618
R1059 vss.n22 vss.n21 0.25832
R1060 vss.n555 vss.n554 0.248562
R1061 vss.n67 vss.n55 0.223756
R1062 vss.n188 vss 0.193102
R1063 vss.n187 vss 0.18715
R1064 vss.n499 vss.n113 0.181206
R1065 vss.n604 vss.n25 0.1605
R1066 vss.n575 vss.n40 0.12599
R1067 vss.n336 vss.n96 0.0491692
R1068 vss.n507 vss.n506 0.0306176
R1069 vss.n348 vss.n262 0.0248346
R1070 vss.n266 vss.n263 0.0248346
R1071 vss.n343 vss.n268 0.0248346
R1072 vss.n297 vss.n296 0.0248346
R1073 vss.n292 vss.n276 0.0248346
R1074 vss.n284 vss.n280 0.0248346
R1075 vss.n446 vss.n445 0.0248346
R1076 vss.n450 vss.n157 0.0248346
R1077 vss.n454 vss.n159 0.0248346
R1078 vss.n500 vss.n499 0.0155588
R1079 vss.n116 vss.n115 0.0155588
R1080 vss.n494 vss.n118 0.0155588
R1081 vss.n493 vss.n119 0.0155588
R1082 vss.n489 vss.n488 0.0155588
R1083 vss.n137 vss.n136 0.0155588
R1084 vss.n483 vss.n139 0.0155588
R1085 vss.n482 vss.n140 0.0155588
R1086 vss.n478 vss.n477 0.0155588
R1087 a_495_638.t1 a_495_638.t0 228.215
R1088 ena.n0 ena.t3 194.3
R1089 ena.n2 ena.t1 62.0385
R1090 ena.n4 ena.t2 5.80898
R1091 ena.n1 ena.t0 4.94781
R1092 ena.n3 ena.t4 4.66216
R1093 ena.n5 ena.n4 1.76704
R1094 ena.n3 ena.n2 1.52716
R1095 ena.n5 ena.n3 1.14731
R1096 ena.n0 ena 0.471358
R1097 ena.n4 ena 0.207161
R1098 ena ena.n5 0.207161
R1099 ena.n2 ena.n1 0.173703
R1100 ena.n1 ena.n0 0.0795843
R1101 a_764_n1158.n0 a_764_n1158.t0 85.9138
R1102 a_764_n1158.n0 a_764_n1158.t2 84.7724
R1103 a_764_n1158.t1 a_764_n1158.n0 84.1936
R1104 XQ_BR1.Emitter.n20 XQ_BR1.Emitter.n19 640.25
R1105 XQ_BR1.Emitter.n7 XQ_BR1.Emitter.t3 228.282
R1106 XQ_BR1.Emitter.n8 XQ_BR1.Emitter.t2 228.22
R1107 XQ_BR1.Emitter.n9 XQ_BR1.Emitter.t0 228.219
R1108 XQ_BR1.Emitter.n10 XQ_BR1.Emitter.t1 228.219
R1109 XQ_BR1.Emitter.n11 XQ_BR1.Emitter.t4 228.215
R1110 XQ_BR1.Emitter.n20 XQ_BR1.Emitter.n14 83.7933
R1111 XQ_BR1.Emitter.n21 XQ_BR1.Emitter.n4 83.5719
R1112 XQ_BR1.Emitter.n22 XQ_BR1.Emitter.n0 83.5719
R1113 XQ_BR1.Emitter.n24 XQ_BR1.Emitter.n23 83.5719
R1114 XQ_BR1.Emitter.n26 XQ_BR1.Emitter.n25 83.5719
R1115 XQ_BR1.Emitter.n25 XQ_BR1.Emitter.n17 73.3165
R1116 XQ_BR1.Emitter.n25 XQ_BR1.Emitter.n24 26.074
R1117 XQ_BR1.Emitter.n22 XQ_BR1.Emitter.n21 26.074
R1118 XQ_BR1.Emitter.n21 XQ_BR1.Emitter.n20 26.074
R1119 XQ_BR1.Emitter.t5 XQ_BR1.Emitter.n22 25.7843
R1120 XQ_BR1.Emitter.n14 XQ_BR1.Emitter.n3 9.3005
R1121 XQ_BR1.Emitter.n32 XQ_BR1.Emitter.n3 9.3005
R1122 XQ_BR1.Emitter.n15 XQ_BR1.Emitter.n3 9.3005
R1123 XQ_BR1.Emitter.n14 XQ_BR1.Emitter.n5 9.3005
R1124 XQ_BR1.Emitter.n32 XQ_BR1.Emitter.n5 9.3005
R1125 XQ_BR1.Emitter.n15 XQ_BR1.Emitter.n5 9.3005
R1126 XQ_BR1.Emitter.n29 XQ_BR1.Emitter.n5 9.3005
R1127 XQ_BR1.Emitter.n14 XQ_BR1.Emitter.n2 9.3005
R1128 XQ_BR1.Emitter.n32 XQ_BR1.Emitter.n2 9.3005
R1129 XQ_BR1.Emitter.n15 XQ_BR1.Emitter.n2 9.3005
R1130 XQ_BR1.Emitter.n29 XQ_BR1.Emitter.n2 9.3005
R1131 XQ_BR1.Emitter.n28 XQ_BR1.Emitter.n14 9.3005
R1132 XQ_BR1.Emitter.n28 XQ_BR1.Emitter.n15 9.3005
R1133 XQ_BR1.Emitter.n29 XQ_BR1.Emitter.n28 9.3005
R1134 XQ_BR1.Emitter.n18 XQ_BR1.Emitter.n14 9.3005
R1135 XQ_BR1.Emitter.n18 XQ_BR1.Emitter.n15 9.3005
R1136 XQ_BR1.Emitter.n18 XQ_BR1.Emitter.n13 9.3005
R1137 XQ_BR1.Emitter.n29 XQ_BR1.Emitter.n18 9.3005
R1138 XQ_BR1.Emitter.n31 XQ_BR1.Emitter.n14 9.3005
R1139 XQ_BR1.Emitter.n32 XQ_BR1.Emitter.n31 9.3005
R1140 XQ_BR1.Emitter.n31 XQ_BR1.Emitter.n15 9.3005
R1141 XQ_BR1.Emitter.n31 XQ_BR1.Emitter.n13 9.3005
R1142 XQ_BR1.Emitter.n6 XQ_BR1.Emitter.t6 5.01718
R1143 XQ_BR1.Emitter.n30 XQ_BR1.Emitter.n29 4.64471
R1144 XQ_BR1.Emitter.n13 XQ_BR1.Emitter.n12 4.64471
R1145 XQ_BR1.Emitter.n27 XQ_BR1.Emitter.n13 4.64471
R1146 XQ_BR1.Emitter.n32 XQ_BR1.Emitter.n1 4.64471
R1147 XQ_BR1.Emitter.n17 XQ_BR1.Emitter.n16 2.24293
R1148 XQ_BR1.Emitter.n14 XQ_BR1.Emitter.n4 1.43912
R1149 XQ_BR1.Emitter.n29 XQ_BR1.Emitter.n17 1.19225
R1150 XQ_BR1.Emitter.n7 XQ_BR1.Emitter.n6 1.08946
R1151 XQ_BR1.Emitter.n23 XQ_BR1.Emitter.n15 1.07024
R1152 XQ_BR1.Emitter.n29 XQ_BR1.Emitter.n26 0.959578
R1153 XQ_BR1.Emitter.n26 XQ_BR1.Emitter.n13 0.885803
R1154 XQ_BR1.Emitter.n23 XQ_BR1.Emitter.n13 0.77514
R1155 XQ_BR1.Emitter XQ_BR1.Emitter.n32 0.756696
R1156 XQ_BR1.Emitter.n15 XQ_BR1.Emitter.n0 0.590702
R1157 XQ_BR1.Emitter XQ_BR1.Emitter.n0 0.498483
R1158 XQ_BR1.Emitter.n32 XQ_BR1.Emitter.n4 0.406264
R1159 XQ_BR1.Emitter.n31 XQ_BR1.Emitter.n11 0.307897
R1160 XQ_BR1.Emitter.n24 XQ_BR1.Emitter.t5 0.290206
R1161 XQ_BR1.Emitter.n10 XQ_BR1.Emitter.n9 0.162265
R1162 XQ_BR1.Emitter.n11 XQ_BR1.Emitter.n10 0.160059
R1163 XQ_BR1.Emitter.n9 XQ_BR1.Emitter.n8 0.158588
R1164 XQ_BR1.Emitter.n8 XQ_BR1.Emitter.n7 0.0990294
R1165 XQ_BR1.Emitter.n6 XQ_BR1.Emitter 0.0239981
R1166 XQ_BR1.Emitter.n16 XQ_BR1.Emitter.n2 0.016881
R1167 XQ_BR1.Emitter.n30 XQ_BR1.Emitter.n3 0.0135838
R1168 XQ_BR1.Emitter.n12 XQ_BR1.Emitter.n5 0.0135838
R1169 XQ_BR1.Emitter.n28 XQ_BR1.Emitter.n27 0.0135838
R1170 XQ_BR1.Emitter.n18 XQ_BR1.Emitter.n1 0.0135838
R1171 XQ_BR1.Emitter.n12 XQ_BR1.Emitter.n3 0.0135838
R1172 XQ_BR1.Emitter.n27 XQ_BR1.Emitter.n2 0.0135838
R1173 XQ_BR1.Emitter.n28 XQ_BR1.Emitter.n1 0.0135838
R1174 XQ_BR1.Emitter.n31 XQ_BR1.Emitter.n30 0.0135838
R1175 XQ_BR1.Emitter.n16 XQ_BR1.Emitter.n5 0.00932056
R1176 vbe1_out vbe1_out.t2 228.484
R1177 vbe1_out.n1 vbe1_out.t3 194.3
R1178 vbe1_out.n0 vbe1_out.t1 83.763
R1179 vbe1_out.n0 vbe1_out.t0 5.02615
R1180 vbe1_out.n1 vbe1_out 0.398938
R1181 vbe1_out.n2 vbe1_out.n0 0.297471
R1182 vbe1_out.n2 vbe1_out.n1 0.124899
R1183 vbe1_out vbe1_out.n2 0.058098
R1184 a_2471_n2640.t0 a_2471_n2640.t1 169.231
R1185 vbe2_out.n1 vbe2_out.t0 228.488
R1186 vbe2_out.n2 vbe2_out.t3 194.535
R1187 vbe2_out.n0 vbe2_out.t2 83.7614
R1188 vbe2_out.n0 vbe2_out.t1 5.03265
R1189 vbe2_out.n1 vbe2_out.n0 0.297705
R1190 vbe2_out vbe2_out.n2 0.107977
R1191 vbe2_out.n2 vbe2_out 0.107977
R1192 vbe2_out vbe2_out.n1 0.041588
R1193 x2.input.n27 x2.input.t0 228.518
R1194 x2.input.n17 x2.input.n14 83.7933
R1195 x2.input.n18 x2.input.n4 83.5719
R1196 x2.input.n19 x2.input.n0 83.5719
R1197 x2.input.n21 x2.input.n20 83.5719
R1198 x2.input.n23 x2.input.n22 83.5719
R1199 x2.input.n24 x2.input.n23 73.3165
R1200 x2.input.n23 x2.input.n21 26.074
R1201 x2.input.n19 x2.input.n18 26.074
R1202 x2.input.n18 x2.input.n17 26.074
R1203 x2.input.t1 x2.input.n19 25.7843
R1204 x2.input.n17 x2.input.n16 20.5696
R1205 x2.input.n14 x2.input.n3 9.3005
R1206 x2.input.n28 x2.input.n3 9.3005
R1207 x2.input.n13 x2.input.n3 9.3005
R1208 x2.input.n15 x2.input.n3 9.3005
R1209 x2.input.n14 x2.input.n7 9.3005
R1210 x2.input.n28 x2.input.n7 9.3005
R1211 x2.input.n13 x2.input.n7 9.3005
R1212 x2.input.n15 x2.input.n7 9.3005
R1213 x2.input.n25 x2.input.n7 9.3005
R1214 x2.input.n14 x2.input.n2 9.3005
R1215 x2.input.n28 x2.input.n2 9.3005
R1216 x2.input.n13 x2.input.n2 9.3005
R1217 x2.input.n15 x2.input.n2 9.3005
R1218 x2.input.n25 x2.input.n2 9.3005
R1219 x2.input.n14 x2.input.n8 9.3005
R1220 x2.input.n28 x2.input.n8 9.3005
R1221 x2.input.n15 x2.input.n8 9.3005
R1222 x2.input.n25 x2.input.n8 9.3005
R1223 x2.input.n14 x2.input.n1 9.3005
R1224 x2.input.n28 x2.input.n1 9.3005
R1225 x2.input.n15 x2.input.n1 9.3005
R1226 x2.input.n11 x2.input.n1 9.3005
R1227 x2.input.n25 x2.input.n1 9.3005
R1228 x2.input.n27 x2.input.n14 9.3005
R1229 x2.input.n28 x2.input.n27 9.3005
R1230 x2.input.n27 x2.input.n13 9.3005
R1231 x2.input.n27 x2.input.n15 9.3005
R1232 x2.input.n27 x2.input.n11 9.3005
R1233 x2.input.n5 x2.input.t2 5.01788
R1234 x2.input.n26 x2.input.n25 4.64593
R1235 x2.input.n11 x2.input.n9 4.64593
R1236 x2.input.n11 x2.input.n10 4.64593
R1237 x2.input.n13 x2.input.n12 4.64593
R1238 x2.input.n6 x2.input.n5 2.03579
R1239 x2.input.n14 x2.input.n4 1.43912
R1240 x2.input.n24 x2.input.n11 1.19225
R1241 x2.input.n20 x2.input.n13 1.07024
R1242 x2.input.n22 x2.input.n11 0.959578
R1243 x2.input.n22 x2.input.n15 0.885803
R1244 x2.input.n20 x2.input.n15 0.77514
R1245 x2.input x2.input.n28 0.756696
R1246 x2.input.n25 x2.input.n24 0.647417
R1247 x2.input.n13 x2.input.n0 0.590702
R1248 x2.input x2.input.n0 0.498483
R1249 x2.input.n28 x2.input.n4 0.406264
R1250 x2.input.n21 x2.input.t1 0.290206
R1251 x2.input.n5 x2.input 0.0236132
R1252 x2.input.n6 x2.input.n2 0.0118636
R1253 x2.input.n26 x2.input.n3 0.011135
R1254 x2.input.n9 x2.input.n7 0.011135
R1255 x2.input.n10 x2.input.n8 0.011135
R1256 x2.input.n12 x2.input.n1 0.011135
R1257 x2.input.n9 x2.input.n3 0.011135
R1258 x2.input.n10 x2.input.n2 0.011135
R1259 x2.input.n12 x2.input.n8 0.011135
R1260 x2.input.n27 x2.input.n26 0.011135
R1261 x2.input.n7 x2.input.n6 0.00942857
R1262 vbg.n0 vbg.t0 194.3
R1263 vbg.n0 vbg.t1 60.3054
R1264 vbg vbg.n0 0.326966
R1265 a_506_n1158.t2 a_506_n1158.n2 228.218
R1266 a_506_n1158.n1 a_506_n1158.t1 120.278
R1267 a_506_n1158.t1 a_506_n1158.n0 120.209
R1268 a_506_n1158.n1 a_506_n1158.t0 85.2046
R1269 a_506_n1158.n0 a_506_n1158.t3 61.8039
R1270 a_506_n1158.n2 a_506_n1158.n0 0.0614063
R1271 a_506_n1158.n2 a_506_n1158.n1 0.0057735
C0 vbg vss 1.96f
C1 vbg ena 0.207f
C2 vss x2.input 8.29f
C3 a_1660_n393# x2.input 0.861f
C4 vbe1_out vss 7.05f
C5 ena x2.input 0.95f
C6 vbe1_out ena 0.256f
C7 a_1537_2302# vss 1.95f
C8 vss XQ_BR1.Emitter 11f
C9 XQ_BR1.Emitter a_1660_n393# 1.75f
C10 a_1537_2302# ena 0.397f
C11 ena XQ_BR1.Emitter 1.32f
C12 a_1537_2302# vbe2_out 0.387f
C13 vss a_1660_n393# 10.5f
C14 vss ena 31.4f
C15 ena a_1660_n393# 1.2f
C16 vss vbe2_out 5.45f
C17 vbe1_out VSUBS 2.24f
C18 vbg VSUBS 0.238f
C19 vbe2_out VSUBS 1.83f
C20 ena VSUBS 7.52f
C21 vss VSUBS 0.192p
C22 x2.input VSUBS 1.21f
C23 a_1660_n393# VSUBS 1.83f
C24 XQ_BR1.Emitter VSUBS 1.33f
C25 a_1537_2302# VSUBS 0.15f
C26 a_506_n1158.t3 VSUBS 0.522f
C27 a_506_n1158.n0 VSUBS 3.19f
C28 a_506_n1158.t1 VSUBS 0.477f
C29 a_506_n1158.n1 VSUBS 0.978f
C30 a_506_n1158.n2 VSUBS 0.172f
C31 x2.input.n1 VSUBS 0.114f
C32 x2.input.n3 VSUBS 0.118f
C33 x2.input.t2 VSUBS 1.21f
C34 x2.input.n5 VSUBS 2.43f
C35 x2.input.n6 VSUBS 1.44f
C36 x2.input.n8 VSUBS 0.118f
C37 x2.input.n14 VSUBS 0.172f
C38 x2.input.n17 VSUBS 0.105f
C39 x2.input.n18 VSUBS 0.118f
C40 x2.input.n19 VSUBS 0.117f
C41 x2.input.n23 VSUBS 0.267f
C42 x2.input.n24 VSUBS 0.122f
C43 x2.input.n25 VSUBS 0.215f
C44 x2.input.n27 VSUBS 0.797f
C45 vbe2_out.t1 VSUBS 1.94f
C46 vbe2_out.n0 VSUBS 2.62f
C47 vbe2_out.n1 VSUBS 0.384f
C48 vbe2_out.n2 VSUBS 0.215f
C49 a_2471_n2640.t1 VSUBS 1.35f
C50 a_2471_n2640.t0 VSUBS 1.35f
C51 vbe1_out.t0 VSUBS 2.39f
C52 vbe1_out.n0 VSUBS 3.21f
C53 vbe1_out.n1 VSUBS 0.374f
C54 vbe1_out.n2 VSUBS 0.3f
C55 XQ_BR1.Emitter.n2 VSUBS 0.106f
C56 XQ_BR1.Emitter.n3 VSUBS 0.129f
C57 XQ_BR1.Emitter.t6 VSUBS 1.63f
C58 XQ_BR1.Emitter.n6 VSUBS 2.68f
C59 XQ_BR1.Emitter.n7 VSUBS 0.718f
C60 XQ_BR1.Emitter.n8 VSUBS 0.371f
C61 XQ_BR1.Emitter.n9 VSUBS 0.447f
C62 XQ_BR1.Emitter.n10 VSUBS 0.449f
C63 XQ_BR1.Emitter.n11 VSUBS 0.626f
C64 XQ_BR1.Emitter.n14 VSUBS 0.232f
C65 XQ_BR1.Emitter.n16 VSUBS 0.393f
C66 XQ_BR1.Emitter.n17 VSUBS 0.376f
C67 XQ_BR1.Emitter.n18 VSUBS 0.148f
C68 XQ_BR1.Emitter.n19 VSUBS -1.82f
C69 XQ_BR1.Emitter.n20 VSUBS 2.03f
C70 XQ_BR1.Emitter.n21 VSUBS 0.159f
C71 XQ_BR1.Emitter.n22 VSUBS 0.158f
C72 XQ_BR1.Emitter.n25 VSUBS 0.36f
C73 XQ_BR1.Emitter.n28 VSUBS 0.129f
C74 XQ_BR1.Emitter.n29 VSUBS 0.118f
C75 XQ_BR1.Emitter.n31 VSUBS 0.495f
C76 a_764_n1158.t0 VSUBS 0.109f
C77 a_764_n1158.n0 VSUBS 4.61f
C78 ena.t0 VSUBS 2.17f
C79 ena.n0 VSUBS 0.678f
C80 ena.n1 VSUBS 3.33f
C81 ena.t1 VSUBS 0.252f
C82 ena.n2 VSUBS 3.62f
C83 ena.t4 VSUBS 2.03f
C84 ena.n3 VSUBS 3.25f
C85 ena.t2 VSUBS 2.62f
C86 ena.n4 VSUBS 7.31f
C87 ena.n5 VSUBS 4.75f
C88 a_495_638.t0 VSUBS 10.6f
C89 vss.n7 VSUBS 2.13f
C90 vss.n8 VSUBS 1.16f
C91 vss.t38 VSUBS 1.94f
C92 vss.n11 VSUBS 1.42f
C93 vss.n13 VSUBS 0.584f
C94 vss.n16 VSUBS 1.83f
C95 vss.t40 VSUBS 1.83f
C96 vss.n20 VSUBS 0.424f
C97 vss.n22 VSUBS 0.131f
C98 vss.n23 VSUBS 0.313f
C99 vss.n24 VSUBS 0.323f
C100 vss.n29 VSUBS 1.83f
C101 vss.n33 VSUBS 1.91f
C102 vss.n34 VSUBS 0.398f
C103 vss.n35 VSUBS 0.899f
C104 vss.n41 VSUBS 0.959f
C105 vss.n42 VSUBS 0.363f
C106 vss.n43 VSUBS 0.689f
C107 vss.n46 VSUBS 0.393f
C108 vss.n48 VSUBS 0.43f
C109 vss.t25 VSUBS 0.326f
C110 vss.n49 VSUBS 0.46f
C111 vss.t9 VSUBS 0.375f
C112 vss.n60 VSUBS 4.49f
C113 vss.n63 VSUBS 1.01f
C114 vss.n64 VSUBS 2.36f
C115 vss.n67 VSUBS 0.263f
C116 vss.n69 VSUBS 0.584f
C117 vss.n72 VSUBS 0.196f
C118 vss.t28 VSUBS -0.149f
C119 vss.n74 VSUBS 0.154f
C120 vss.n76 VSUBS 0.426f
C121 vss.n77 VSUBS 0.146f
C122 vss.n78 VSUBS 0.229f
C123 vss.n79 VSUBS 0.222f
C124 vss.n80 VSUBS 2.06f
C125 vss.t10 VSUBS 0.534f
C126 vss.n87 VSUBS 0.301f
C127 vss.n89 VSUBS 0.18f
C128 vss.n91 VSUBS 0.212f
C129 vss.n92 VSUBS 0.146f
C130 vss.t37 VSUBS 2.81f
C131 vss.t36 VSUBS 1.94f
C132 vss.n124 VSUBS 1.86f
C133 vss.n125 VSUBS 1.28f
C134 vss.n126 VSUBS 0.705f
C135 vss.n127 VSUBS 0.205f
C136 vss.n130 VSUBS 0.492f
C137 vss.n133 VSUBS 0.108f
C138 vss.n134 VSUBS 0.123f
C139 vss.n148 VSUBS 0.116f
C140 vss.t34 VSUBS 1.94f
C141 vss.n178 VSUBS 0.326f
C142 vss.n186 VSUBS 0.376f
C143 vss.n187 VSUBS 3.21f
C144 vss.n188 VSUBS 2.36f
C145 vss.n189 VSUBS 0.378f
C146 vss.n194 VSUBS 0.301f
C147 vss.n200 VSUBS 0.301f
C148 vss.n201 VSUBS 0.301f
C149 vss.n207 VSUBS 0.301f
C150 vss.n208 VSUBS 0.222f
C151 vss.t35 VSUBS 0.268f
C152 vss.n390 VSUBS 0.301f
C153 vss.t5 VSUBS 0.196f
C154 vss.n399 VSUBS 0.231f
C155 vss.n400 VSUBS 0.301f
C156 vss.n406 VSUBS 0.301f
C157 vss.n407 VSUBS 0.301f
C158 vss.n408 VSUBS 0.229f
C159 vss.n411 VSUBS 0.475f
C160 vss.n412 VSUBS 0.486f
C161 vss.n415 VSUBS 0.475f
C162 vss.n416 VSUBS 3.13f
C163 vss.n507 VSUBS 0.155f
C164 vss.n529 VSUBS 0.585f
C165 vss.n530 VSUBS 0.45f
C166 vss.n536 VSUBS 0.301f
C167 vss.n537 VSUBS 0.301f
C168 vss.n538 VSUBS 0.301f
C169 vss.n545 VSUBS 0.301f
C170 vss.n546 VSUBS 0.301f
C171 vss.n550 VSUBS 0.134f
C172 vss.n551 VSUBS 0.299f
C173 vss.n552 VSUBS 0.313f
C174 vss.n553 VSUBS 0.318f
C175 vss.n555 VSUBS 0.785f
C176 vss.n557 VSUBS 0.686f
C177 vss.t39 VSUBS -1.41f
C178 vss.n558 VSUBS 0.167f
C179 vss.n562 VSUBS 0.115f
C180 vss.n563 VSUBS 0.15f
C181 vss.n566 VSUBS 0.1f
C182 vss.n571 VSUBS 0.88f
C183 vss.t32 VSUBS 2.61f
C184 vss.n573 VSUBS 0.127f
C185 vss.t41 VSUBS 0.568f
C186 vss.n581 VSUBS 0.407f
C187 vss.n582 VSUBS 0.111f
C188 vss.t6 VSUBS 0.136f
C189 vss.n586 VSUBS 0.375f
C190 vss.n590 VSUBS 0.101f
C191 vss.n592 VSUBS 0.646f
C192 vss.n593 VSUBS 0.288f
C193 vss.n595 VSUBS 0.507f
C194 vss.n598 VSUBS 0.114f
C195 vss.n601 VSUBS 4.39f
C196 vss.n602 VSUBS 1.69f
C197 vss.n603 VSUBS 1.62f
C198 vss.t4 VSUBS 0.414f
C199 vss.n613 VSUBS 0.221f
C200 vss.n615 VSUBS 0.483f
C201 vss.n616 VSUBS 0.12f
C202 vss.n617 VSUBS 0.232f
C203 vss.t23 VSUBS 1.83f
C204 vss.n619 VSUBS 1.83f
C205 vss.n622 VSUBS 0.1f
C206 vss.n624 VSUBS 0.117f
C207 vss.n626 VSUBS 2.18f
C208 vss.n627 VSUBS 3.91f
C209 vss.n628 VSUBS 1.6f
C210 vss.n629 VSUBS 0.63f
C211 a_1429_n4304.t1 VSUBS 11.6f
.ends

*testbanch circuit
V1 vdd GND 1.8
V2 vbg GND 1.2
x1 vdd vbe1 vdd vbg vbe2 GND tempsensor_rcx

*simulation def 
.func mu(vbe1,vbe2) = 10.7906/(10.7906+vbe1/(vbe2-vbe1))
.func T(mu) = 714.015*mu-259.802
.control
option TEMP=25
op
let ttrim = T(mu(V(vbe1),V(vbe2)))-25
*** DEBUG - search for linear mode trasistor
*set altshow
*show > /tmp/tras.txt

dc temp -40 125 10
plot V(vbe1) V(vbe2)-V(vbe1) V(vbe1)+10.7906*(V(vbe2)-V(vbe1))
plot T(mu(V(vbe1),V(vbe2)))-op1.ttrim
plot T(mu(V(vbe1),V(vbe2)))-\"temp-sweep\"-op1.ttrim
plot V(vbe1) V(vbe2)


.endc