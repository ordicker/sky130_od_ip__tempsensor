magic
tech sky130A
magscale 1 2
timestamp 1713170137
<< locali >>
rect 4838 2878 9524 3150
rect 3510 2824 10034 2878
rect 3510 2700 3594 2824
rect 9964 2700 10034 2824
rect 3510 2524 10034 2700
rect 3514 2432 10034 2524
rect 3514 2430 6604 2432
rect 3514 1864 3680 2430
rect 4134 2276 4560 2430
rect 4022 2272 4560 2276
rect 4022 2096 4674 2272
rect 4134 2092 4674 2096
rect 5014 2268 5474 2430
rect 5938 2270 6604 2430
rect 7066 2372 10034 2432
rect 4134 1856 4560 2092
rect 5014 2088 5596 2268
rect 5014 1860 5474 2088
rect 5938 2084 6724 2270
rect 5938 1878 6604 2084
rect 7066 1886 7684 2372
rect 7844 2270 8022 2372
rect 8280 2274 8458 2372
rect 8718 2274 8896 2372
rect 9152 2272 9330 2372
rect 9588 2268 9766 2372
rect 9930 1878 10034 2372
rect 5938 1864 6072 1878
rect 9370 1678 10036 1680
rect 3520 1570 6484 1666
rect 3520 1096 3674 1570
rect 4134 1096 5480 1570
rect 5930 1096 6484 1570
rect 3520 1034 6484 1096
rect 3520 892 3674 1034
rect 3520 760 3794 892
rect 3522 706 3794 760
rect 3522 568 3674 706
rect 5930 582 6484 1034
rect 7304 582 8418 1672
rect 9232 582 10036 1678
rect 5930 568 10038 582
rect 3522 326 10038 568
rect 3522 324 10034 326
rect 3526 228 10034 324
rect 3526 104 3616 228
rect 9906 104 10034 228
rect 3526 62 10034 104
rect 4402 -40 9102 62
<< viali >>
rect 3594 2700 9964 2824
rect 3616 104 9906 228
<< metal1 >>
rect 8418 5050 8428 5254
rect 9338 5050 9348 5254
rect 8362 4670 8372 4938
rect 9282 4670 9292 4938
rect 4848 3794 5048 3994
rect 8934 3810 8944 3986
rect 9136 3810 9146 3986
rect 3564 2852 3764 2862
rect 3550 2826 10004 2852
rect 3550 2824 5960 2826
rect 6280 2824 10004 2826
rect 3550 2700 3594 2824
rect 9964 2700 10004 2824
rect 3550 2698 5960 2700
rect 6280 2698 10004 2700
rect 3550 2672 10004 2698
rect 3564 2662 3764 2672
rect 3876 2556 5756 2570
rect 3876 2476 5758 2556
rect 3876 2364 3956 2476
rect 3584 2270 3796 2272
rect 3874 2270 3956 2364
rect 5664 2360 5758 2476
rect 3584 2226 3956 2270
rect 3584 2096 3952 2226
rect 3584 2094 3796 2096
rect 3584 1402 3656 2094
rect 3874 2004 3952 2096
rect 4736 2040 4840 2358
rect 4900 2092 5122 2270
rect 5662 2196 5758 2360
rect 5934 2444 7564 2588
rect 5934 2270 6056 2444
rect 6748 2326 6920 2444
rect 3808 1608 4008 1860
rect 4680 1842 4888 2040
rect 3582 1226 3794 1402
rect 3834 1142 3980 1608
rect 4680 1514 4712 1842
rect 4858 1514 4888 1842
rect 5028 1832 5120 2092
rect 5662 2000 5756 2196
rect 5820 2092 6056 2270
rect 5934 1832 6056 2092
rect 6788 2002 6878 2326
rect 7100 2274 7232 2276
rect 6944 2098 7232 2274
rect 7396 2214 7562 2444
rect 7396 2108 9858 2214
rect 7100 1878 7232 2098
rect 5028 1682 6056 1832
rect 5028 1680 5120 1682
rect 4680 1484 4888 1514
rect 4022 1228 5596 1400
rect 4656 1092 4846 1228
rect 5654 1146 5766 1682
rect 5934 1656 6056 1682
rect 6546 1864 7232 1878
rect 5934 1400 6002 1656
rect 6546 1642 6568 1864
rect 7198 1642 7232 1864
rect 7840 1876 8022 2058
rect 8282 1876 8464 2060
rect 8718 1876 8900 2056
rect 9152 1876 9334 2054
rect 9586 1876 9768 2056
rect 7840 1868 9768 1876
rect 7840 1752 8526 1868
rect 7842 1708 8526 1752
rect 5818 1226 6004 1400
rect 5944 1092 6008 1094
rect 4656 1038 6008 1092
rect 4656 1036 4846 1038
rect 4002 636 5542 966
rect 5944 888 6008 1038
rect 5820 712 6010 888
rect 5944 710 6008 712
rect 6546 664 7232 1642
rect 8502 1646 8526 1708
rect 9156 1750 9768 1868
rect 9156 1708 9766 1750
rect 9156 1646 9188 1708
rect 8502 662 9188 1646
rect 4326 602 5068 636
rect 4326 350 4744 602
rect 5042 350 5068 602
rect 4326 326 5068 350
rect 3580 262 3780 286
rect 3580 256 9976 262
rect 3580 244 9980 256
rect 3580 228 7746 244
rect 8172 228 9980 244
rect 3580 104 3616 228
rect 9906 104 9980 228
rect 3580 84 9978 104
rect 7942 -332 7952 -86
rect 8844 -332 8854 -86
rect 4398 -1558 4598 -1358
rect 8482 -1556 8492 -1344
rect 8690 -1556 8700 -1344
rect 5944 -2356 5954 -2228
rect 6274 -2356 6284 -2228
<< via1 >>
rect 8428 5050 9338 5254
rect 8372 4670 9282 4938
rect 8944 3810 9136 3986
rect 5960 2824 6280 2826
rect 5960 2700 6280 2824
rect 5960 2698 6280 2700
rect 4712 1514 4858 1842
rect 6568 1642 7198 1864
rect 8526 1646 9156 1868
rect 4744 350 5042 602
rect 7746 228 8172 244
rect 7746 110 8172 228
rect 7952 -332 8844 -86
rect 8492 -1556 8690 -1344
rect 5954 -2356 6274 -2228
<< metal2 >>
rect 5090 5254 9500 5278
rect 5090 5050 8428 5254
rect 9338 5050 9500 5254
rect 5090 5020 9500 5050
rect 5090 3210 5396 5020
rect 8372 4938 9282 4948
rect 8372 4660 9282 4670
rect 8380 4584 9280 4660
rect 7748 4580 9280 4584
rect 7746 4292 9280 4580
rect 7746 4282 9256 4292
rect 7316 3210 7608 3216
rect 5090 2956 7608 3210
rect 5090 1864 5396 2956
rect 5960 2834 6280 2836
rect 5956 2826 6284 2834
rect 5956 2698 5960 2826
rect 6280 2698 6284 2826
rect 4706 1842 5414 1864
rect 4706 1514 4712 1842
rect 4858 1514 5414 1842
rect 4706 1506 5414 1514
rect 4712 1504 4968 1506
rect 4744 616 4968 1504
rect 4744 602 5042 616
rect 4744 340 5042 350
rect 5956 -2218 6284 2698
rect 6568 1864 7198 1874
rect 6568 1632 7198 1642
rect 6936 -1344 7190 1632
rect 7316 -78 7608 2956
rect 7746 244 8186 4282
rect 8944 3992 9136 3996
rect 8944 3986 9138 3992
rect 9136 3810 9138 3986
rect 8944 1878 9138 3810
rect 8526 1868 9156 1878
rect 8526 1636 9156 1646
rect 8172 110 8186 244
rect 7746 100 8172 110
rect 7952 -78 8844 -76
rect 7316 -86 9074 -78
rect 7316 -332 7952 -86
rect 8844 -332 9074 -86
rect 7316 -352 9074 -332
rect 8492 -1344 8690 -1334
rect 6934 -1556 8492 -1344
rect 8690 -1556 8694 -1344
rect 6934 -1560 8694 -1556
rect 8492 -1566 8690 -1560
rect 5954 -2228 6284 -2218
rect 6274 -2352 6284 -2228
rect 5954 -2366 6274 -2356
use buffer  x1
timestamp 1713093572
transform -1 0 9832 0 -1 -1930
box 726 -1956 5440 496
use buffer  x2
timestamp 1713093572
transform -1 0 10280 0 -1 3412
box 726 -1956 5440 496
use sky130_fd_pr__pfet_01v8_lvt_3VR9VM  XM1
timestamp 1713031642
transform 1 0 6834 0 1 2179
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_lvt_6VRZAW  XM2
timestamp 1713031642
transform 0 1 8807 -1 0 2160
box -296 -1191 296 1191
use sky130_fd_pr__pfet_01v8_3HMWVM  XM3
timestamp 1713031642
transform 1 0 4788 0 1 2179
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_69TQ3K  XM4
timestamp 1713031642
transform 1 0 3908 0 1 1314
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_69TQ3K  XM5
timestamp 1713031642
transform 1 0 5706 0 1 1316
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_NXBWHY  XM6
timestamp 1713031642
transform 1 0 4808 0 1 798
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM7
timestamp 1713031642
transform 1 0 5708 0 1 2179
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_3HMWVM  XM8
timestamp 1713031642
transform 1 0 3910 0 1 2183
box -296 -319 296 319
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ_BL1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1698934549
transform 1 0 6224 0 1 330
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ_BR1
timestamp 1698934549
transform 1 0 8160 0 1 310
box 0 0 1340 1340
<< labels >>
flabel metal1 3808 1660 4008 1860 0 FreeSans 256 0 0 0 vbg
port 5 nsew
flabel metal1 4516 332 4716 532 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal1 3580 86 3780 286 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 3564 2662 3764 2862 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 4398 -1558 4598 -1358 0 FreeSans 256 0 0 0 Vbe1
port 3 nsew
flabel metal1 4848 3794 5048 3994 0 FreeSans 256 0 0 0 Vbe2
port 2 nsew
<< end >>
