magic
tech sky130A
magscale 1 2
timestamp 1713856378
<< nwell >>
rect -584 2916 6610 3202
rect -584 -4744 -298 2916
rect 6324 -4744 6610 2916
rect -584 -5030 6610 -4744
<< nsubdiff >>
rect -547 3145 6573 3165
rect -547 3111 -467 3145
rect 6493 3111 6573 3145
rect -547 3091 6573 3111
rect -547 3085 -473 3091
rect -547 -4913 -527 3085
rect -493 -4913 -473 3085
rect -547 -4919 -473 -4913
rect 6499 3085 6573 3091
rect 6499 -4913 6519 3085
rect 6553 -4913 6573 3085
rect 6499 -4919 6573 -4913
rect -547 -4939 6573 -4919
rect -547 -4973 -467 -4939
rect 6493 -4973 6573 -4939
rect -547 -4993 6573 -4973
<< nsubdiffcont >>
rect -467 3111 6493 3145
rect -527 -4913 -493 3085
rect 6519 -4913 6553 3085
rect -467 -4973 6493 -4939
<< locali >>
rect -527 3111 -467 3145
rect 6493 3111 6553 3145
rect -527 3085 -493 3111
rect 6519 3085 6553 3111
rect 496 2712 600 2716
rect -50 2662 600 2712
rect -50 2130 6 2662
rect -50 1678 404 2130
rect 5228 1822 5966 2062
rect 234 1374 404 1678
rect 5226 1668 5966 1822
rect 5230 534 5440 1668
rect 5878 1512 5966 1668
rect 5774 1342 5966 1512
rect 5878 1074 5966 1342
rect 5770 904 5966 1074
rect 5878 644 5966 904
rect 302 38 5440 534
rect 5774 474 5966 644
rect 5878 200 5966 474
rect 320 -50 5440 38
rect 5770 30 5966 200
rect 320 -602 448 -50
rect 888 -200 1344 -50
rect 1784 -200 2240 -50
rect 2684 -74 5440 -50
rect 778 -382 1450 -200
rect 888 -388 1450 -382
rect 1784 -382 2346 -200
rect 888 -602 1344 -388
rect 1784 -594 2240 -382
rect 2684 -612 4102 -74
rect 4542 -222 5440 -74
rect 4432 -386 5440 -222
rect 5878 -234 5966 30
rect 4542 -606 5440 -386
rect 5774 -404 5966 -234
rect 4542 -612 5438 -606
rect 5878 -630 5966 -404
rect 370 -1288 472 -744
rect 876 -1288 2240 -748
rect 2686 -1288 3536 -746
rect 370 -1554 3536 -1288
rect 370 -1692 472 -1554
rect 370 -1874 554 -1692
rect 370 -2022 472 -1874
rect 2686 -2022 3536 -1554
rect 4356 -2022 4858 -732
rect 5694 -2022 5942 -760
rect 370 -2238 5942 -2022
rect 370 -2248 5940 -2238
rect 370 -2250 472 -2248
rect 664 -2834 1020 -2248
rect 664 -2882 1332 -2834
rect 812 -3292 1332 -2882
rect 812 -3532 1342 -3292
rect 812 -3816 940 -3532
rect 300 -4660 1278 -4346
rect -527 -4939 -493 -4913
rect 6519 -4939 6553 -4913
rect -527 -4973 -467 -4939
rect 6493 -4973 6553 -4939
<< viali >>
rect 6 2130 1216 2662
<< metal1 >>
rect -36 2662 1274 2704
rect -36 2130 6 2662
rect 1216 2130 1274 2662
rect 3850 2362 3860 2594
rect 4722 2362 4732 2594
rect -36 2080 1274 2130
rect 3842 2026 3852 2288
rect 4758 2026 4768 2288
rect 70 1368 174 1604
rect 5594 1586 5714 1612
rect -64 1154 550 1368
rect 4090 1148 4100 1366
rect 4596 1148 4606 1366
rect 5124 1346 5556 1518
rect 5112 1156 5122 1346
rect 5394 1332 5556 1346
rect 5394 1156 5464 1332
rect 5124 1076 5464 1156
rect 5124 890 5556 1076
rect 5124 646 5464 890
rect 1790 326 1800 504
rect 2538 326 2548 504
rect 5124 460 5554 646
rect 5124 206 5464 460
rect 564 -14 2530 144
rect 5124 20 5556 206
rect 564 -20 710 -14
rect 566 -98 710 -20
rect 520 -202 710 -98
rect 420 -224 710 -202
rect 420 -380 708 -224
rect 422 -964 478 -380
rect 520 -478 708 -380
rect 1492 -442 1614 -114
rect 1668 -386 1990 -204
rect 2402 -208 2528 -14
rect 2712 -162 3038 -120
rect 4262 -128 4378 -124
rect 2712 -198 2760 -162
rect 1466 -658 1644 -442
rect 1848 -616 1990 -386
rect 2404 -476 2524 -208
rect 2572 -378 2760 -198
rect 2684 -552 2760 -378
rect 2986 -552 3038 -162
rect 4252 -156 4392 -128
rect 2684 -602 3038 -552
rect 3776 -400 4200 -214
rect 2684 -616 3030 -602
rect 1456 -852 1466 -658
rect 1636 -852 1646 -658
rect 1848 -746 3030 -616
rect 1850 -750 3030 -746
rect 1466 -864 1644 -852
rect 422 -1140 552 -964
rect 610 -1196 706 -886
rect 1558 -960 2348 -958
rect 772 -1142 2348 -960
rect 2432 -962 2608 -868
rect 2684 -962 3030 -750
rect 2432 -1122 3030 -962
rect 3776 -1118 4128 -400
rect 4252 -466 4268 -156
rect 4368 -466 4392 -156
rect 4252 -486 4392 -466
rect 5124 -228 5464 20
rect 5124 -414 5550 -228
rect 5124 -1092 5464 -414
rect 5594 -452 5610 1586
rect 5706 -452 5716 1586
rect 5594 -500 5716 -452
rect 5594 -502 5714 -500
rect 2432 -1126 2740 -1122
rect 2432 -1136 2716 -1126
rect 772 -1144 1596 -1142
rect 576 -1224 706 -1196
rect 366 -1402 708 -1224
rect 1348 -1358 1596 -1144
rect 2432 -1230 2608 -1136
rect 3632 -1156 4248 -1118
rect 2676 -1358 2762 -1356
rect 366 -2252 472 -1402
rect 1344 -1478 2762 -1358
rect 824 -1954 2278 -1610
rect 2676 -1692 2762 -1478
rect 2578 -1862 2762 -1692
rect 3632 -1706 3678 -1156
rect 4204 -1706 4248 -1156
rect 3632 -1728 4248 -1706
rect 3776 -1738 4128 -1728
rect 4968 -1752 5610 -1092
rect 2578 -1870 2756 -1862
rect 954 -2124 1240 -1954
rect 952 -2232 1240 -2124
rect 952 -2238 1242 -2232
rect 1716 -2238 3192 -2178
rect 366 -2412 602 -2252
rect 952 -2254 3192 -2238
rect 366 -2546 472 -2412
rect 952 -2526 1138 -2254
rect 1904 -2304 3192 -2254
rect 1904 -2526 1994 -2304
rect 2854 -2360 3192 -2304
rect 2860 -2434 3192 -2360
rect 952 -2544 1994 -2526
rect 364 -2788 578 -2546
rect 952 -2548 1242 -2544
rect 952 -2994 1238 -2548
rect 4772 -2902 4782 -2648
rect 5658 -2902 5668 -2648
rect 5672 -2884 5942 -2688
rect 350 -3236 1238 -2994
rect 350 -3242 1164 -3236
rect 328 -3592 578 -3580
rect 328 -3800 1444 -3592
rect 5006 -3788 5016 -3580
rect 5526 -3788 5536 -3580
rect 328 -3822 578 -3800
rect 302 -4454 620 -4404
rect 302 -4622 1356 -4454
rect 302 -4624 1340 -4622
rect 2062 -4630 2072 -4452
rect 2810 -4630 2820 -4452
<< via1 >>
rect 3860 2362 4722 2594
rect 3852 2026 4758 2288
rect 4100 1148 4596 1366
rect 5122 1156 5394 1346
rect 1800 326 2538 504
rect 2760 -552 2986 -162
rect 1466 -852 1636 -658
rect 4268 -466 4368 -156
rect 5610 -452 5706 1586
rect 3678 -1706 4204 -1156
rect 1138 -2526 1904 -2254
rect 4794 -2566 5656 -2334
rect 4782 -2902 5658 -2648
rect 5016 -3788 5526 -3580
rect 2072 -4630 2810 -4452
<< metal2 >>
rect 4394 2620 4954 2630
rect 3860 2594 4394 2614
rect 4722 2362 4954 2366
rect 3860 2356 4954 2362
rect 3860 2352 4722 2356
rect 3852 2288 4758 2298
rect 4758 2274 4760 2284
rect 3852 2010 4760 2020
rect 5610 1586 5708 1608
rect 4100 1368 4596 1376
rect 4100 1366 5392 1368
rect 4596 1356 5392 1366
rect 4596 1346 5394 1356
rect 4596 1156 5122 1346
rect 4596 1148 5394 1156
rect 4100 1146 5394 1148
rect 4100 1144 5392 1146
rect 4100 1138 4596 1144
rect 1800 504 2538 514
rect 1800 316 2538 326
rect 1426 -658 1660 -640
rect 1426 -852 1466 -658
rect 1636 -852 1660 -658
rect 1426 -2244 1660 -852
rect 1806 -1432 2534 316
rect 2760 -156 2986 -152
rect 4268 -156 5610 -146
rect 2758 -162 4268 -156
rect 2758 -478 2760 -162
rect 2986 -466 4268 -162
rect 4368 -452 5610 -156
rect 5706 -452 5708 1586
rect 4368 -466 5708 -452
rect 2986 -478 4368 -466
rect 5610 -470 5708 -466
rect 2760 -562 2986 -552
rect 3678 -1156 4204 -1146
rect 1806 -1490 2782 -1432
rect 1806 -1700 2780 -1490
rect 1138 -2254 1904 -2244
rect 1138 -2536 1904 -2526
rect 2068 -4442 2780 -1700
rect 3678 -1716 4204 -1706
rect 3808 -3578 4064 -1716
rect 4780 -2334 5950 -2302
rect 4780 -2564 4794 -2334
rect 5656 -2556 5950 -2334
rect 4794 -2576 5656 -2566
rect 4782 -2638 5164 -2632
rect 4782 -2642 5658 -2638
rect 5164 -2648 5658 -2642
rect 4782 -2912 5658 -2902
rect 5016 -3578 5526 -3570
rect 3808 -3580 5526 -3578
rect 3808 -3772 5016 -3580
rect 3808 -3780 4064 -3772
rect 5016 -3798 5526 -3788
rect 2068 -4452 2810 -4442
rect 2068 -4630 2072 -4452
rect 2068 -4640 2810 -4630
rect 2068 -4642 2780 -4640
<< via2 >>
rect 4394 2594 4954 2620
rect 4394 2366 4722 2594
rect 4722 2366 4954 2594
rect 3852 2026 4758 2274
rect 4758 2026 4760 2274
rect 3852 2020 4760 2026
rect 5310 -2554 5646 -2336
rect 4782 -2648 5164 -2642
rect 4782 -2902 5164 -2648
<< metal3 >>
rect 4384 2620 4964 2625
rect 4384 2366 4394 2620
rect 4954 2588 4964 2620
rect 4954 2366 5652 2588
rect 4384 2361 5652 2366
rect 4400 2360 5652 2361
rect 3842 2274 4770 2279
rect 3832 2020 3852 2274
rect 4760 2020 5144 2274
rect 3832 1994 5144 2020
rect 4772 -2637 5144 1994
rect 5310 -2331 5652 2360
rect 5300 -2336 5656 -2331
rect 5300 -2554 5310 -2336
rect 5646 -2554 5656 -2336
rect 5300 -2559 5656 -2554
rect 5310 -2570 5652 -2559
rect 4772 -2642 5174 -2637
rect 4772 -2902 4782 -2642
rect 5164 -2902 5174 -2642
rect 4772 -2907 5174 -2902
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0
timestamp 1713474431
transform 1 0 553 0 1 -2341
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_1
timestamp 1713474431
transform 1 0 1133 0 1 -2725
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_2
timestamp 1713474431
transform 1 0 1033 0 1 -3639
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_3
timestamp 1713474431
transform 1 0 129 0 1 1563
box -183 -183 183 183
use buffer  x1
timestamp 1713290077
transform -1 0 5736 0 -1 780
box 726 -1956 5440 496
use buffer  x2
timestamp 1713290077
transform -1 0 6670 0 -1 -4162
box 726 -1956 5440 496
use sky130_fd_pr__pfet_01v8_lvt_3VR9VM  XM11
timestamp 1713290077
transform 1 0 4320 0 1 -307
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_lvt_6VRZAW  XM22
timestamp 1713290077
transform 1 0 5662 0 1 551
box -296 -1191 296 1191
use sky130_fd_pr__pfet_01v8_3HMWVM  XM33
timestamp 1713290077
transform 1 0 1560 0 1 -293
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_69TQ3K  XM44
timestamp 1713290077
transform 1 0 664 0 1 -1058
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_69TQ3K  XM55
timestamp 1713290077
transform 1 0 2460 0 1 -1054
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_QXBCRM  XM66
timestamp 1713290077
transform 1 0 1568 0 1 -1784
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM77
timestamp 1713290077
transform 1 0 2460 0 1 -291
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_3HMWVM  XM88
timestamp 1713290077
transform 1 0 672 0 1 -293
box -296 -319 296 319
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ_BL1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1698934549
transform 1 0 3272 0 1 -2100
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ_BR1
timestamp 1698934549
transform 1 0 4616 0 1 -2100
box 0 0 1340 1340
<< labels >>
flabel metal1 302 -4604 502 -4404 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 370 -2770 570 -2570 0 FreeSans 256 0 0 0 vbg
port 5 nsew
flabel metal1 356 -3218 556 -3018 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal1 336 -3806 536 -3606 0 FreeSans 256 0 0 0 vbe1_out
port 3 nsew
flabel metal1 -62 1158 138 1358 0 FreeSans 256 0 0 0 vbe2_out
port 2 nsew
flabel locali 30 2508 230 2708 0 FreeSans 256 0 0 0 vss
port 1 nsew
<< end >>
