magic
tech sky130A
magscale 1 2
timestamp 1713031642
<< nwell >>
rect -296 -1191 296 1191
<< pmoslvt >>
rect -100 772 100 972
rect -100 336 100 536
rect -100 -100 100 100
rect -100 -536 100 -336
rect -100 -972 100 -772
<< pdiff >>
rect -158 960 -100 972
rect -158 784 -146 960
rect -112 784 -100 960
rect -158 772 -100 784
rect 100 960 158 972
rect 100 784 112 960
rect 146 784 158 960
rect 100 772 158 784
rect -158 524 -100 536
rect -158 348 -146 524
rect -112 348 -100 524
rect -158 336 -100 348
rect 100 524 158 536
rect 100 348 112 524
rect 146 348 158 524
rect 100 336 158 348
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
rect -158 -348 -100 -336
rect -158 -524 -146 -348
rect -112 -524 -100 -348
rect -158 -536 -100 -524
rect 100 -348 158 -336
rect 100 -524 112 -348
rect 146 -524 158 -348
rect 100 -536 158 -524
rect -158 -784 -100 -772
rect -158 -960 -146 -784
rect -112 -960 -100 -784
rect -158 -972 -100 -960
rect 100 -784 158 -772
rect 100 -960 112 -784
rect 146 -960 158 -784
rect 100 -972 158 -960
<< pdiffc >>
rect -146 784 -112 960
rect 112 784 146 960
rect -146 348 -112 524
rect 112 348 146 524
rect -146 -88 -112 88
rect 112 -88 146 88
rect -146 -524 -112 -348
rect 112 -524 146 -348
rect -146 -960 -112 -784
rect 112 -960 146 -784
<< nsubdiff >>
rect -260 1121 -164 1155
rect 164 1121 260 1155
rect -260 1059 -226 1121
rect 226 1059 260 1121
rect -260 -1121 -226 -1059
rect 226 -1121 260 -1059
rect -260 -1155 -164 -1121
rect 164 -1155 260 -1121
<< nsubdiffcont >>
rect -164 1121 164 1155
rect -260 -1059 -226 1059
rect 226 -1059 260 1059
rect -164 -1155 164 -1121
<< poly >>
rect -100 1053 100 1069
rect -100 1019 -84 1053
rect 84 1019 100 1053
rect -100 972 100 1019
rect -100 725 100 772
rect -100 691 -84 725
rect 84 691 100 725
rect -100 675 100 691
rect -100 617 100 633
rect -100 583 -84 617
rect 84 583 100 617
rect -100 536 100 583
rect -100 289 100 336
rect -100 255 -84 289
rect 84 255 100 289
rect -100 239 100 255
rect -100 181 100 197
rect -100 147 -84 181
rect 84 147 100 181
rect -100 100 100 147
rect -100 -147 100 -100
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect -100 -197 100 -181
rect -100 -255 100 -239
rect -100 -289 -84 -255
rect 84 -289 100 -255
rect -100 -336 100 -289
rect -100 -583 100 -536
rect -100 -617 -84 -583
rect 84 -617 100 -583
rect -100 -633 100 -617
rect -100 -691 100 -675
rect -100 -725 -84 -691
rect 84 -725 100 -691
rect -100 -772 100 -725
rect -100 -1019 100 -972
rect -100 -1053 -84 -1019
rect 84 -1053 100 -1019
rect -100 -1069 100 -1053
<< polycont >>
rect -84 1019 84 1053
rect -84 691 84 725
rect -84 583 84 617
rect -84 255 84 289
rect -84 147 84 181
rect -84 -181 84 -147
rect -84 -289 84 -255
rect -84 -617 84 -583
rect -84 -725 84 -691
rect -84 -1053 84 -1019
<< locali >>
rect -260 1121 -164 1155
rect 164 1121 260 1155
rect -260 1059 -226 1121
rect 226 1059 260 1121
rect -100 1019 -84 1053
rect 84 1019 100 1053
rect -146 960 -112 976
rect -146 768 -112 784
rect 112 960 146 976
rect 112 768 146 784
rect -100 691 -84 725
rect 84 691 100 725
rect -100 583 -84 617
rect 84 583 100 617
rect -146 524 -112 540
rect -146 332 -112 348
rect 112 524 146 540
rect 112 332 146 348
rect -100 255 -84 289
rect 84 255 100 289
rect -100 147 -84 181
rect 84 147 100 181
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect -100 -289 -84 -255
rect 84 -289 100 -255
rect -146 -348 -112 -332
rect -146 -540 -112 -524
rect 112 -348 146 -332
rect 112 -540 146 -524
rect -100 -617 -84 -583
rect 84 -617 100 -583
rect -100 -725 -84 -691
rect 84 -725 100 -691
rect -146 -784 -112 -768
rect -146 -976 -112 -960
rect 112 -784 146 -768
rect 112 -976 146 -960
rect -100 -1053 -84 -1019
rect 84 -1053 100 -1019
rect -260 -1121 -226 -1059
rect 226 -1121 260 -1059
rect -260 -1155 -164 -1121
rect 164 -1155 260 -1121
<< viali >>
rect -84 1019 84 1053
rect -146 784 -112 960
rect 112 784 146 960
rect -84 691 84 725
rect -84 583 84 617
rect -146 348 -112 524
rect 112 348 146 524
rect -84 255 84 289
rect -84 147 84 181
rect -146 -88 -112 88
rect 112 -88 146 88
rect -84 -181 84 -147
rect -84 -289 84 -255
rect -146 -524 -112 -348
rect 112 -524 146 -348
rect -84 -617 84 -583
rect -84 -725 84 -691
rect -146 -960 -112 -784
rect 112 -960 146 -784
rect -84 -1053 84 -1019
<< metal1 >>
rect -96 1053 96 1059
rect -96 1019 -84 1053
rect 84 1019 96 1053
rect -96 1013 96 1019
rect -152 960 -106 972
rect -152 784 -146 960
rect -112 784 -106 960
rect -152 772 -106 784
rect 106 960 152 972
rect 106 784 112 960
rect 146 784 152 960
rect 106 772 152 784
rect -96 725 96 731
rect -96 691 -84 725
rect 84 691 96 725
rect -96 685 96 691
rect -96 617 96 623
rect -96 583 -84 617
rect 84 583 96 617
rect -96 577 96 583
rect -152 524 -106 536
rect -152 348 -146 524
rect -112 348 -106 524
rect -152 336 -106 348
rect 106 524 152 536
rect 106 348 112 524
rect 146 348 152 524
rect 106 336 152 348
rect -96 289 96 295
rect -96 255 -84 289
rect 84 255 96 289
rect -96 249 96 255
rect -96 181 96 187
rect -96 147 -84 181
rect 84 147 96 181
rect -96 141 96 147
rect -152 88 -106 100
rect -152 -88 -146 88
rect -112 -88 -106 88
rect -152 -100 -106 -88
rect 106 88 152 100
rect 106 -88 112 88
rect 146 -88 152 88
rect 106 -100 152 -88
rect -96 -147 96 -141
rect -96 -181 -84 -147
rect 84 -181 96 -147
rect -96 -187 96 -181
rect -96 -255 96 -249
rect -96 -289 -84 -255
rect 84 -289 96 -255
rect -96 -295 96 -289
rect -152 -348 -106 -336
rect -152 -524 -146 -348
rect -112 -524 -106 -348
rect -152 -536 -106 -524
rect 106 -348 152 -336
rect 106 -524 112 -348
rect 146 -524 152 -348
rect 106 -536 152 -524
rect -96 -583 96 -577
rect -96 -617 -84 -583
rect 84 -617 96 -583
rect -96 -623 96 -617
rect -96 -691 96 -685
rect -96 -725 -84 -691
rect 84 -725 96 -691
rect -96 -731 96 -725
rect -152 -784 -106 -772
rect -152 -960 -146 -784
rect -112 -960 -106 -784
rect -152 -972 -106 -960
rect 106 -784 152 -772
rect 106 -960 112 -784
rect 146 -960 152 -784
rect 106 -972 152 -960
rect -96 -1019 96 -1013
rect -96 -1053 -84 -1019
rect 84 -1053 96 -1019
rect -96 -1059 96 -1053
<< properties >>
string FIXED_BBOX -243 -1138 243 1138
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 1.0 l 1.0 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
