* NGSPICE file created from sky130_od_ip__tempsensor_ext_vp.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_QXBCRM a_n1000_n188# a_n1160_n274# a_1000_n100# a_n1058_n100#
X0 a_1000_n100# a_n1000_n188# a_n1058_n100# a_n1160_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
C0 a_1000_n100# a_n1160_n274# 0.177f
C1 a_n1058_n100# a_n1160_n274# 0.177f
C2 a_n1000_n188# a_n1160_n274# 5.78f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_B5H3CA w_n1196_n319# a_n1000_n197# a_1000_n100#
+ a_n1058_n100# VSUBS
X0 a_1000_n100# a_n1000_n197# a_n1058_n100# w_n1196_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
C0 w_n1196_n319# a_n1000_n197# 3.21f
C1 a_n1000_n197# VSUBS 2.69f
C2 w_n1196_n319# VSUBS 5.96f
.ends

.subckt buffer input output vdd vbias vss m1_772_n974#
XXM1 input vss m1_2942_n986# m1_772_n974# sky130_fd_pr__nfet_01v8_QXBCRM
XXM2 output vss output m1_2942_n986# sky130_fd_pr__nfet_01v8_QXBCRM
XXM3 vdd m1_772_n974# vdd m1_772_n974# vss sky130_fd_pr__pfet_01v8_lvt_B5H3CA
XXM4 vdd m1_772_n974# output vdd vss sky130_fd_pr__pfet_01v8_lvt_B5H3CA
XXM5 vbias vss m1_2942_n986# vss sky130_fd_pr__nfet_01v8_QXBCRM
C0 input m1_772_n974# 0.403f
C1 m1_772_n974# vdd 2.09f
C2 vbias input 0.133f
C3 output vdd 0.23f
C4 output m1_2942_n986# 0.337f
C5 vbias m1_2942_n986# 0.348f
C6 output m1_772_n974# 0.363f
C7 vbias vss 8.67f
C8 m1_772_n974# vss 4.96f
C9 vdd vss 12.9f
C10 m1_2942_n986# vss 2.04f
C11 output vss 6.28f
C12 input vss 6.04f
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
C0 Emitter Base 0.897f
C1 Base Collector 1.11f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_6VRZAW a_100_n536# w_n296_n1191# a_n100_675# a_100_336#
+ a_n158_n536# a_n158_772# a_n100_n633# a_n100_239# a_n100_n197# a_100_n100# a_n158_336#
+ a_100_n972# a_n158_n100# a_100_772# a_n158_n972# a_n100_n1069# VSUBS
X0 a_100_336# a_n100_239# a_n158_336# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_772# a_n100_675# a_n158_772# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_n536# a_n100_n633# a_n158_n536# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_100_n972# a_n100_n1069# a_n158_n972# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 w_n296_n1191# a_n100_239# 0.262f
C1 a_n100_n633# a_n100_n1069# 0.205f
C2 a_n100_n633# a_n100_n197# 0.205f
C3 a_n100_n1069# w_n296_n1191# 0.348f
C4 a_n100_n633# w_n296_n1191# 0.262f
C5 a_n100_675# w_n296_n1191# 0.348f
C6 w_n296_n1191# a_n100_n197# 0.262f
C7 a_n100_675# a_n100_239# 0.205f
C8 a_n100_n197# a_n100_239# 0.205f
C9 a_n100_n1069# VSUBS 0.257f
C10 a_n100_n633# VSUBS 0.204f
C11 a_n100_n197# VSUBS 0.204f
C12 a_n100_239# VSUBS 0.204f
C13 a_n100_675# VSUBS 0.257f
C14 w_n296_n1191# VSUBS 5.73f
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_3VR9VM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
+ VSUBS
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 w_n296_n319# a_n100_n197# 0.434f
C1 a_n100_n197# VSUBS 0.311f
C2 w_n296_n319# VSUBS 1.65f
.ends

.subckt sky130_fd_pr__pfet_01v8_3HMWVM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
+ VSUBS
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 w_n296_n319# a_n100_n197# 0.434f
C1 a_n100_n197# VSUBS 0.311f
C2 w_n296_n319# VSUBS 1.65f
.ends

.subckt sky130_fd_pr__nfet_01v8_69TQ3K a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_100_n100# a_n260_n274# 0.146f
C1 a_n158_n100# a_n260_n274# 0.146f
C2 a_n100_n188# a_n260_n274# 0.724f
.ends

.subckt sky130_od_ip__tempsensor_ext_vp vdd vss vbe2_out vbe1_out ena vbg
Xx1 x1/input vbe2_out vdd ena vss x1/m1_772_n974# buffer
Xx2 x2/input vbe1_out vdd ena vss x2/m1_772_n974# buffer
XXQ_BR1 x1/input vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXQ_BL1 x2/input vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXM22 vdd vdd m1_1668_n386# vdd x1/input x1/input m1_1668_n386# m1_1668_n386# m1_1668_n386#
+ vdd x1/input vdd x1/input vdd x1/input m1_1668_n386# vss sky130_fd_pr__pfet_01v8_lvt_6VRZAW
XXM11 vdd m1_1668_n386# vdd x2/input vss sky130_fd_pr__pfet_01v8_lvt_3VR9VM
XXM33 vdd ena m1_1668_n386# vdd vss sky130_fd_pr__pfet_01v8_3HMWVM
XXM44 vss m1_772_n1144# m1_420_n380# vbg sky130_fd_pr__nfet_01v8_69TQ3K
XXM55 vss m1_1668_n386# m1_772_n1144# m1_1668_n386# sky130_fd_pr__nfet_01v8_69TQ3K
XXM66 ena vss m1_772_n1144# vss sky130_fd_pr__nfet_01v8_QXBCRM
XXM77 vdd m1_420_n380# m1_1668_n386# vdd vss sky130_fd_pr__pfet_01v8_3HMWVM
XXM88 vdd m1_420_n380# vdd m1_420_n380# vss sky130_fd_pr__pfet_01v8_3HMWVM
C0 m1_1668_n386# vdd 3.66f
C1 ena m1_420_n380# 0.105f
C2 x2/m1_772_n974# vdd 0.453f
C3 ena m1_772_n1144# 1.17f
C4 ena vbe1_out 0.115f
C5 x1/m1_772_n974# x1/input 0.508f
C6 ena x2/input 0.862f
C7 x1/m1_772_n974# vdd 0.208f
C8 m1_420_n380# vdd 3.31f
C9 vdd m1_772_n1144# 0.296f
C10 ena vbg 0.163f
C11 vbe1_out vdd 0.857f
C12 m1_1668_n386# m1_420_n380# 0.281f
C13 x2/input vdd 0.762f
C14 m1_1668_n386# m1_772_n1144# 0.216f
C15 vbg vdd 0.279f
C16 m1_1668_n386# x2/input 0.834f
C17 ena x1/input 0.187f
C18 ena vdd 2.09f
C19 x2/m1_772_n974# x2/input 0.592f
C20 ena m1_1668_n386# 0.58f
C21 vdd x1/input 2.38f
C22 m1_420_n380# vbg 0.156f
C23 m1_1668_n386# x1/input 1.62f
C24 m1_420_n380# vss 0.988f
C25 vdd vss 42.1f
C26 m1_1668_n386# vss 3.91f
C27 m1_772_n1144# vss 3.26f
C28 vbg vss 2.11f
C29 x1/input vss 5.98f
C30 ena vss 29f
C31 x2/m1_772_n974# vss 4.81f
C32 x2/m1_2942_n986# vss 0.485f
C33 vbe1_out vss 5.85f
C34 x2/input vss 6.58f
C35 x1/m1_772_n974# vss 4.82f
C36 x1/m1_2942_n986# vss 0.497f
C37 vbe2_out vss 5.76f
.ends

