magic
tech sky130A
magscale 1 2
timestamp 1713295635
<< locali >>
rect 5228 1822 5966 2062
rect 5226 1668 5966 1822
rect 5230 534 5440 1668
rect 5878 1512 5966 1668
rect 5774 1342 5966 1512
rect 5878 1074 5966 1342
rect 5770 904 5966 1074
rect 5878 644 5966 904
rect 302 38 5440 534
rect 5774 474 5966 644
rect 5878 200 5966 474
rect 320 -50 5440 38
rect 5770 30 5966 200
rect 320 -602 448 -50
rect 888 -200 1344 -50
rect 1784 -200 2240 -50
rect 2684 -74 5440 -50
rect 778 -382 1450 -200
rect 888 -388 1450 -382
rect 1784 -382 2346 -200
rect 888 -602 1344 -388
rect 1784 -594 2240 -382
rect 2684 -612 4102 -74
rect 4542 -222 5440 -74
rect 4432 -386 5440 -222
rect 5878 -234 5966 30
rect 4542 -606 5440 -386
rect 5774 -404 5966 -234
rect 4542 -612 5438 -606
rect 5878 -630 5966 -404
rect 370 -1288 472 -744
rect 876 -1288 2240 -748
rect 2686 -1288 3536 -746
rect 370 -1554 3536 -1288
rect 370 -1692 472 -1554
rect 370 -1874 554 -1692
rect 370 -2022 472 -1874
rect 2686 -2022 3536 -1554
rect 4356 -2022 4858 -732
rect 5694 -2022 5942 -760
rect 370 -2238 5942 -2022
rect 370 -2248 5940 -2238
rect 370 -2250 472 -2248
rect 300 -4660 1278 -4346
<< metal1 >>
rect 3850 2362 3860 2594
rect 4722 2362 4732 2594
rect 6034 2320 6288 2338
rect 4708 2028 6288 2320
rect 5594 1586 5714 1612
rect -108 1146 506 1360
rect 5124 1332 5556 1518
rect 5124 1076 5464 1332
rect 5124 890 5556 1076
rect 5124 646 5464 890
rect 1298 310 1308 490
rect 2024 310 2034 490
rect 5124 460 5554 646
rect 5124 206 5464 460
rect 564 -14 2530 144
rect 5124 20 5556 206
rect 564 -20 710 -14
rect 566 -98 710 -20
rect 520 -202 710 -98
rect 420 -224 710 -202
rect 420 -380 708 -224
rect 422 -964 478 -380
rect 520 -478 708 -380
rect 1492 -442 1614 -114
rect 1668 -386 1990 -204
rect 2402 -208 2528 -14
rect 2712 -162 3038 -120
rect 4262 -128 4378 -124
rect 2712 -198 2760 -162
rect 1466 -658 1644 -442
rect 1848 -616 1990 -386
rect 2404 -476 2524 -208
rect 2572 -378 2760 -198
rect 2684 -552 2760 -378
rect 2986 -552 3038 -162
rect 4252 -156 4392 -128
rect 2684 -602 3038 -552
rect 3776 -400 4200 -214
rect 2684 -616 3030 -602
rect 1456 -852 1466 -658
rect 1636 -852 1646 -658
rect 1848 -746 3030 -616
rect 1850 -750 3030 -746
rect 1466 -864 1644 -852
rect 422 -1140 552 -964
rect 610 -1196 706 -886
rect 1558 -960 2348 -958
rect 772 -1142 2348 -960
rect 2432 -962 2608 -868
rect 2684 -962 3030 -750
rect 2432 -1122 3030 -962
rect 3776 -1118 4128 -400
rect 4252 -466 4268 -156
rect 4368 -466 4392 -156
rect 4252 -486 4392 -466
rect 5124 -228 5464 20
rect 5124 -414 5550 -228
rect 5124 -1092 5464 -414
rect 5594 -452 5610 1586
rect 5706 -452 5716 1586
rect 5594 -500 5716 -452
rect 5594 -502 5714 -500
rect 2432 -1126 2740 -1122
rect 2432 -1136 2716 -1126
rect 772 -1144 1596 -1142
rect 576 -1298 740 -1196
rect -12 -1440 740 -1298
rect 1348 -1358 1596 -1144
rect 2432 -1230 2608 -1136
rect 2676 -1358 2762 -1356
rect -12 -1446 706 -1440
rect -12 -2722 114 -1446
rect 1344 -1478 2762 -1358
rect 824 -1954 2278 -1610
rect 2676 -1692 2762 -1478
rect 2578 -1862 2762 -1692
rect 3632 -1728 4248 -1118
rect 3776 -1738 4128 -1728
rect 4968 -1752 5610 -1092
rect 2578 -1870 2756 -1862
rect 954 -2232 1240 -1954
rect 342 -2238 1242 -2232
rect 1716 -2238 3192 -2178
rect 342 -2254 3192 -2238
rect 342 -2526 1138 -2254
rect 1904 -2304 3192 -2254
rect 1904 -2526 1994 -2304
rect 2854 -2360 3192 -2304
rect 2860 -2434 3192 -2360
rect 342 -2544 1994 -2526
rect 342 -2548 1242 -2544
rect 4784 -2566 4794 -2334
rect 5656 -2566 5666 -2334
rect 6034 -2688 6288 2028
rect 5672 -2692 6302 -2688
rect -12 -2964 492 -2722
rect 5672 -2884 6304 -2692
rect 6104 -2892 6304 -2884
rect 282 -3592 1442 -3590
rect 278 -3788 1442 -3592
rect 278 -3792 478 -3788
rect 302 -4452 502 -4404
rect 302 -4454 1340 -4452
rect 302 -4618 1304 -4454
rect 2032 -4618 2042 -4454
rect 302 -4624 1340 -4618
<< via1 >>
rect 3860 2362 4722 2594
rect 1308 310 2024 490
rect 2760 -552 2986 -162
rect 1466 -852 1636 -658
rect 4268 -466 4368 -156
rect 5610 -452 5706 1586
rect 1138 -2526 1904 -2254
rect 4794 -2566 5656 -2334
rect 1304 -4618 2032 -4454
<< metal2 >>
rect 3860 2594 6236 2614
rect 4722 2362 6236 2594
rect 3860 2352 4722 2362
rect 5610 1586 5708 1608
rect 740 492 2036 506
rect 736 490 2036 492
rect 736 310 1308 490
rect 2024 486 2036 490
rect 2024 310 2038 486
rect 736 292 2036 310
rect 736 -2788 938 292
rect 2760 -156 2986 -152
rect 4268 -156 5610 -146
rect 2758 -162 4268 -156
rect 2758 -478 2760 -162
rect 2986 -466 4268 -162
rect 4368 -452 5610 -156
rect 5706 -452 5708 1586
rect 4368 -466 5708 -452
rect 2986 -478 4368 -466
rect 5610 -470 5708 -466
rect 2760 -562 2986 -552
rect 1426 -658 1660 -640
rect 1426 -852 1466 -658
rect 1636 -852 1660 -658
rect 1426 -2244 1660 -852
rect 1138 -2254 1904 -2244
rect 5950 -2302 6214 2362
rect 1138 -2536 1904 -2526
rect 4780 -2334 6214 -2302
rect 4780 -2564 4794 -2334
rect 5656 -2556 6214 -2334
rect 5656 -2564 6192 -2556
rect 4794 -2576 5656 -2566
rect 736 -2806 1436 -2788
rect 736 -3120 1440 -2806
rect 1298 -4226 1440 -3120
rect 1298 -4454 2026 -4226
rect 1298 -4618 1304 -4454
rect 2032 -4618 2038 -4454
rect 1298 -4622 2038 -4618
rect 1304 -4626 2038 -4622
rect 1304 -4628 2032 -4626
use buffer  x1
timestamp 1713290077
transform -1 0 5736 0 -1 780
box 726 -1956 5440 496
use buffer  x2
timestamp 1713290077
transform -1 0 6670 0 -1 -4162
box 726 -1956 5440 496
use sky130_fd_pr__pfet_01v8_lvt_3VR9VM  XM11
timestamp 1713290077
transform 1 0 4320 0 1 -307
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_lvt_6VRZAW  XM22
timestamp 1713290077
transform 1 0 5662 0 1 551
box -296 -1191 296 1191
use sky130_fd_pr__pfet_01v8_3HMWVM  XM33
timestamp 1713290077
transform 1 0 1560 0 1 -293
box -296 -319 296 319
use sky130_fd_pr__nfet_01v8_69TQ3K  XM44
timestamp 1713290077
transform 1 0 664 0 1 -1058
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_69TQ3K  XM55
timestamp 1713290077
transform 1 0 2460 0 1 -1054
box -296 -310 296 310
use sky130_fd_pr__nfet_01v8_QXBCRM  XM66
timestamp 1713290077
transform 1 0 1568 0 1 -1784
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_3HMWVM  XM77
timestamp 1713290077
transform 1 0 2460 0 1 -291
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_3HMWVM  XM88
timestamp 1713290077
transform 1 0 672 0 1 -293
box -296 -319 296 319
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ_BL1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1698934549
transform 1 0 3272 0 1 -2100
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  XQ_BR1
timestamp 1698934549
transform 1 0 4616 0 1 -2100
box 0 0 1340 1340
<< labels >>
flabel metal1 302 -4604 502 -4404 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 278 -3792 478 -3592 0 FreeSans 256 0 0 0 Vbe1
port 3 nsew
flabel metal1 -106 1150 94 1350 0 FreeSans 256 0 0 0 Vbe2
port 2 nsew
flabel metal1 6104 -2892 6304 -2692 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 346 -2526 546 -2326 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal1 284 -2946 484 -2746 0 FreeSans 256 0 0 0 vbg
port 5 nsew
<< end >>
